
-- 
-- Definition of  FC_controller
-- 
--      Sat May 11 15:31:53 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity FC_controller is
   port (
      clk : IN std_logic ;
      rst : IN std_logic ;
      initiate : INOUT std_logic ;
      enable_read : OUT std_logic ;
      address_out : INOUT std_logic_vector (15 DOWNTO 0) ;
      data_in : IN std_logic_vector (255 DOWNTO 0) ;
      answer : OUT std_logic_vector (3 DOWNTO 0) ;
      done_comp : INOUT std_logic ;
      cnn_address : IN std_logic_vector (15 DOWNTO 0)) ;
end FC_controller ;

architecture a_FC_controller of FC_controller is
   signal enable_read_EXMPLR, answer_3_EXMPLR, answer_2_EXMPLR, 
      answer_1_EXMPLR, answer_0_EXMPLR, max_calc_start, start_comp, state_0, 
      nx18145, state_2, nx18146, nx4, sub_state_2, num_out_2, sub_state_0, 
      nx18153, nx20, nx36, nx50, nx68, num_in_2, nx86, alu_sel, nx18155, 
      nx98, nx104, ready_signal, nx18158, nx122, nx132, 
      enable_decoder_dst_booth, output_17, output_16, output_15, output_14, 
      output_13, output_12, output_11, output_10, output_9, output_8, 
      output_7, output_6, output_5, output_4, output_3, output_2, output_1, 
      output_0, nx246, alu_inp1_0, address_in_0, nx18159, nx284, nx294, 
      nx306, nx326, nx336, nx338, neuron_address_0, nx360, nx362, temp_0, 
      nx388, num_out_0, num_in_0, nx406, nx420, alu_inp2_0, nx442, 
      alu_inp1_1, address_in_1, neuron_address_1, nx18161, nx444, temp_1, 
      nx468, num_out_1, num_in_1, nx500, alu_inp1_2, address_in_2, 
      neuron_address_2, nx18162, nx516, temp_2, nx538, nx554, nx570, 
      num_out_3, num_in_3, nx596, alu_inp1_3, address_in_3, neuron_address_3, 
      nx18163, temp_3, nx620, nx636, nx644, num_out_4, num_in_4, alu_inp1_4, 
      address_in_4, neuron_address_4, nx18165, nx670, temp_4, nx692, nx708, 
      nx724, nx742, num_out_5, num_in_5, nx748, alu_inp1_5, address_in_5, 
      neuron_address_5, nx18167, temp_5, nx772, nx788, nx796, num_out_6, 
      num_in_6, alu_inp1_6, address_in_6, neuron_address_6, nx18169, nx822, 
      temp_6, nx844, nx860, nx876, num_out_7, num_in_7, nx898, alu_inp1_7, 
      address_in_7, neuron_address_7, nx18171, temp_7, nx922, nx938, nx946, 
      num_out_8, num_in_8, alu_inp1_8, address_in_8, neuron_address_8, 
      nx18173, nx972, temp_8, nx994, nx1010, nx1026, nx1044, num_out_9, 
      num_in_9, nx1052, alu_inp1_9, address_in_9, neuron_address_9, nx18175, 
      temp_9, nx1076, nx1092, nx1100, num_out_10, num_in_10, alu_inp1_10, 
      address_in_10, neuron_address_10, nx18177, nx1126, temp_10, nx1148, 
      nx1164, nx1180, num_out_11, num_in_11, nx1202, alu_inp1_11, 
      address_in_11, neuron_address_11, nx18178, temp_11, nx1226, nx1242, 
      nx1250, num_out_12, num_in_12, alu_inp1_12, address_in_12, 
      neuron_address_12, nx18179, nx1276, temp_12, nx1298, nx1314, nx1330, 
      nx1348, num_out_13, num_in_13, nx1354, alu_inp1_13, address_in_13, 
      neuron_address_13, nx18180, temp_13, nx1378, nx1394, nx1402, 
      num_out_14, num_in_14, alu_inp1_14, address_in_14, neuron_address_14, 
      nx18181, nx1428, temp_14, nx1450, nx1466, nx1482, num_out_15, 
      num_in_15, nx1504, alu_inp1_15, address_in_15, neuron_address_15, 
      nx18182, temp_15, nx1528, nx1544, nx1576, nx1582, nx1592, nx1602, 
      nx1612, nx1672, nx1678, nx1714, max_calc_answer_0, max_calc_state_1, 
      max_calc_state_0, max_calc_state_2, nx18183, nx18187, nx1758, nx18189, 
      nx18191, nx1774, nx1782, max_calc_comparator_first_inp1_0, 
      label_1_output_0, sel_dst_0, nx1860, label_1_input_0, 
      booth_booth_integration_output_0_12, 
      booth_booth_integrtaion_0_shift_reg_output_9, 
      booth_booth_integrtaion_0_shift_Reg_count_9, output_8_dup_12688, 
      booth_booth_integrtaion_0_shift_Reg_count_8, output_7_dup_12689, 
      booth_booth_integrtaion_0_shift_Reg_count_7, output_6_dup_12690, 
      booth_booth_integrtaion_0_shift_Reg_count_6, output_5_dup_12691, 
      booth_booth_integrtaion_0_shift_Reg_count_5, output_4_dup_12692, 
      booth_booth_integrtaion_0_shift_Reg_count_4, output_3_dup_12693, 
      booth_booth_integrtaion_0_shift_Reg_count_3, output_2_dup_12694, 
      booth_booth_integrtaion_0_shift_Reg_count_2, output_1_dup_12695, 
      booth_booth_integrtaion_0_shift_Reg_count_1, 
      booth_booth_integrtaion_0_shift_reg_output_0, 
      booth_booth_integrtaion_0_shift_Reg_count_0, 
      booth_booth_integration_output_0_13, 
      booth_booth_integration_output_0_14, 
      booth_booth_integration_output_0_15, 
      booth_booth_integration_output_0_16, booth_output_0, booth_output_1, 
      booth_output_2, booth_output_3, booth_output_4, booth_output_5, 
      booth_output_6, booth_output_7, booth_output_8, booth_output_9, 
      booth_output_10, booth_output_11, neuron_11, nx1980, neuron_10, nx1998, 
      neuron_9, nx2016, neuron_8, nx2034, neuron_7, nx2052, neuron_6, nx2070, 
      neuron_5, nx2088, neuron_4, nx2106, neuron_3, nx2124, neuron_2, nx2142, 
      neuron_1, nx2160, neuron_0, nx2178, nx2204, 
      booth_booth_integration_output_0_17, nx18195, nx2212, nx2218, nx2228, 
      booth_booth_integration_output_0_18, nx18196, nx2238, nx2242, nx2256, 
      booth_booth_integration_output_0_19, nx18197, nx2266, nx2276, 
      booth_booth_integration_output_0_20, nx18198, nx2286, nx2304, 
      booth_booth_integration_output_0_21, nx18199, nx2310, nx2314, nx2324, 
      booth_booth_integration_output_0_22, nx18200, nx2334, nx2352, 
      booth_booth_integration_output_0_23, nx18201, nx2358, nx2362, nx2372, 
      booth_booth_integration_output_0_24, nx18203, nx2382, nx2400, 
      booth_booth_integration_output_0_25, nx18205, nx2406, nx2410, nx2420, 
      booth_booth_integration_output_0_26, nx18207, nx2430, nx2448, 
      booth_booth_integration_output_0_27, nx18209, nx2454, nx2458, nx2468, 
      booth_output_28, nx18210, nx2478, nx2496, booth_output_29, nx18211, 
      nx2502, nx2506, nx2516, nx18212, nx2526, nx2544, nx2552, nx2556, 
      nx2568, nx2584, nx2592, nx2608, nx2616, nx2632, nx2640, nx2656, nx2664, 
      nx2680, nx2688, nx2700, nx2712, nx2728, nx2734, nx2740, neuron_15, 
      neuron_14, nx2770, neuron_13, nx2788, neuron_12, nx2806, nx2818, 
      label_1_input_state_machine_0, nx2830, max_calc_ans1_0, nx2862, 
      nx18213, nx2876, max_calc_ans6_0, max_calc_ans5_0, 
      max_calc_comparator_fifth_inp1_0, label_9_output_0, label_9_input_0, 
      booth_booth_integration_output_8_12, 
      booth_booth_integrtaion_8_shift_reg_output_9, 
      booth_booth_integrtaion_8_shift_Reg_count_9, output_8_dup_12912, 
      booth_booth_integrtaion_8_shift_Reg_count_8, output_7_dup_12913, 
      booth_booth_integrtaion_8_shift_Reg_count_7, output_6_dup_12914, 
      booth_booth_integrtaion_8_shift_Reg_count_6, output_5_dup_12915, 
      booth_booth_integrtaion_8_shift_Reg_count_5, output_4_dup_12916, 
      booth_booth_integrtaion_8_shift_Reg_count_4, output_3_dup_12917, 
      booth_booth_integrtaion_8_shift_Reg_count_3, output_2_dup_12918, 
      booth_booth_integrtaion_8_shift_Reg_count_2, output_1_dup_12919, 
      booth_booth_integrtaion_8_shift_Reg_count_1, 
      booth_booth_integrtaion_8_shift_reg_output_0, 
      booth_booth_integrtaion_8_shift_Reg_count_0, 
      booth_booth_integration_output_8_13, 
      booth_booth_integration_output_8_14, 
      booth_booth_integration_output_8_15, 
      booth_booth_integration_output_8_16, booth_output_0_dup_12263, 
      booth_output_1_dup_12262, booth_output_2_dup_12261, 
      booth_output_3_dup_12260, booth_output_4_dup_12259, 
      booth_output_5_dup_12258, booth_output_6_dup_12257, 
      booth_output_7_dup_12256, booth_output_8_dup_12255, 
      booth_output_9_dup_12254, booth_output_10_dup_12253, 
      booth_output_11_dup_12252, nx2988, nx3000, nx3012, nx3024, nx3036, 
      nx3048, nx3060, nx3072, nx3084, nx3096, nx3108, nx3120, nx3146, 
      booth_booth_integration_output_8_17, nx18215, nx3154, nx3160, nx3170, 
      booth_booth_integration_output_8_18, nx18217, nx3180, nx3184, nx3198, 
      booth_booth_integration_output_8_19, nx18219, nx3208, nx3218, 
      booth_booth_integration_output_8_20, nx18221, nx3228, nx3246, 
      booth_booth_integration_output_8_21, nx18223, nx3252, nx3256, nx3266, 
      booth_booth_integration_output_8_22, nx18225, nx3276, nx3294, 
      booth_booth_integration_output_8_23, nx18227, nx3300, nx3304, nx3314, 
      booth_booth_integration_output_8_24, nx18228, nx3324, nx3342, 
      booth_booth_integration_output_8_25, nx18229, nx3348, nx3352, nx3362, 
      booth_booth_integration_output_8_26, nx18230, nx3372, nx3390, 
      booth_booth_integration_output_8_27, nx18231, nx3396, nx3400, nx3410, 
      booth_output_28_dup_12251, nx18232, nx3420, nx3438, 
      booth_output_29_dup_12250, nx18233, nx3444, nx3448, nx3458, nx18235, 
      nx3468, nx3486, nx3494, nx3498, nx3510, nx3526, nx3534, nx3550, nx3558, 
      nx3574, nx3582, nx3598, nx3606, nx3622, nx3630, nx3642, nx3654, nx3670, 
      nx3676, nx3682, nx3700, nx3712, nx3724, nx3736, 
      label_9_input_state_machine_0, nx3748, label_10_output_14, 
      label_10_input_14, label_10_input_state_machine_14, label_10_output_0, 
      label_10_input_0, booth_booth_integration_output_9_12, 
      booth_booth_integrtaion_9_shift_reg_output_9, 
      booth_booth_integrtaion_9_shift_Reg_count_9, output_8_dup_12940, 
      booth_booth_integrtaion_9_shift_Reg_count_8, output_7_dup_12941, 
      booth_booth_integrtaion_9_shift_Reg_count_7, output_6_dup_12942, 
      booth_booth_integrtaion_9_shift_Reg_count_6, output_5_dup_12943, 
      booth_booth_integrtaion_9_shift_Reg_count_5, output_4_dup_12944, 
      booth_booth_integrtaion_9_shift_Reg_count_4, output_3_dup_12945, 
      booth_booth_integrtaion_9_shift_Reg_count_3, output_2_dup_12946, 
      booth_booth_integrtaion_9_shift_Reg_count_2, output_1_dup_12947, 
      booth_booth_integrtaion_9_shift_Reg_count_1, 
      booth_booth_integrtaion_9_shift_reg_output_0, 
      booth_booth_integrtaion_9_shift_Reg_count_0, 
      booth_booth_integration_output_9_13, 
      booth_booth_integration_output_9_14, 
      booth_booth_integration_output_9_15, 
      booth_booth_integration_output_9_16, booth_output_0_dup_12282, 
      booth_output_1_dup_12281, booth_output_2_dup_12280, 
      booth_output_3_dup_12279, booth_output_4_dup_12278, 
      booth_output_5_dup_12277, booth_output_6_dup_12276, 
      booth_output_7_dup_12275, booth_output_8_dup_12274, 
      booth_output_9_dup_12273, booth_output_10_dup_12272, 
      booth_output_11_dup_12271, nx3868, nx3880, nx3892, nx3904, nx3916, 
      nx3928, nx3940, nx3952, nx3964, nx3976, nx3988, nx4000, nx4026, 
      booth_booth_integration_output_9_17, nx18239, nx4034, nx4040, nx4050, 
      booth_booth_integration_output_9_18, nx18241, nx4060, nx4064, nx4078, 
      booth_booth_integration_output_9_19, nx18242, nx4088, nx4098, 
      booth_booth_integration_output_9_20, nx18243, nx4108, nx4126, 
      booth_booth_integration_output_9_21, nx18244, nx4132, nx4136, nx4146, 
      booth_booth_integration_output_9_22, nx18245, nx4156, nx4174, 
      booth_booth_integration_output_9_23, nx18246, nx4180, nx4184, nx4194, 
      booth_booth_integration_output_9_24, nx18247, nx4204, nx4222, 
      booth_booth_integration_output_9_25, nx18249, nx4228, nx4232, nx4242, 
      booth_booth_integration_output_9_26, nx18251, nx4252, nx4270, 
      booth_booth_integration_output_9_27, nx18253, nx4276, nx4280, nx4290, 
      booth_output_28_dup_12270, nx18254, nx4300, nx4318, 
      booth_output_29_dup_12269, nx18255, nx4324, nx4328, nx4338, nx18256, 
      nx4348, nx4366, nx4374, nx4378, nx4390, nx4406, nx4414, nx4430, nx4438, 
      nx4454, nx4462, nx4478, nx4486, nx4502, nx4510, nx4522, nx4534, nx4550, 
      nx4556, nx4562, nx4580, nx4592, nx4604, nx4614, 
      label_10_input_state_machine_0, nx4626, label_10_output_1, 
      label_10_input_1, label_10_input_state_machine_1, nx4648, nx4652, 
      nx4670, label_10_output_2, label_10_input_2, 
      label_10_input_state_machine_2, nx18259, nx4680, nx4684, 
      label_10_output_3, label_10_input_3, label_10_input_state_machine_3, 
      nx4712, nx4716, nx4734, label_10_output_4, label_10_input_4, 
      label_10_input_state_machine_4, nx18261, nx4744, nx4748, 
      label_10_output_5, label_10_input_5, label_10_input_state_machine_5, 
      nx4776, nx4780, nx4798, label_10_output_6, label_10_input_6, 
      label_10_input_state_machine_6, nx18264, nx4808, nx4812, 
      label_10_output_7, label_10_input_7, label_10_input_state_machine_7, 
      nx4840, nx4844, nx4862, label_10_output_8, label_10_input_8, 
      label_10_input_state_machine_8, nx18266, nx4872, nx4876, 
      label_10_output_9, label_10_input_9, label_10_input_state_machine_9, 
      nx4904, nx4908, nx4926, label_10_output_10, label_10_input_10, 
      label_10_input_state_machine_10, nx18268, nx4936, nx4940, 
      label_10_output_11, label_10_input_11, label_10_input_state_machine_11, 
      nx4968, nx4972, nx4990, label_10_output_12, label_10_input_12, 
      label_10_input_state_machine_12, nx18271, nx5000, nx5004, 
      label_10_output_13, label_10_input_13, label_10_input_state_machine_13, 
      nx5032, nx5036, nx5054, nx5056, nx5058, nx5062, 
      max_calc_comparator_fifth_inp1_14, label_9_output_14, label_9_input_14, 
      label_9_input_state_machine_14, label_9_output_1, label_9_input_1, 
      label_9_input_state_machine_1, nx5098, nx5102, nx5120, 
      label_9_output_2, label_9_input_2, label_9_input_state_machine_2, 
      nx18277, nx5130, nx5134, label_9_output_3, label_9_input_3, 
      label_9_input_state_machine_3, nx5162, nx5166, nx5184, 
      label_9_output_4, label_9_input_4, label_9_input_state_machine_4, 
      nx18280, nx5194, nx5198, label_9_output_5, label_9_input_5, 
      label_9_input_state_machine_5, nx5226, nx5230, nx5248, 
      label_9_output_6, label_9_input_6, label_9_input_state_machine_6, 
      nx18282, nx5258, nx5262, label_9_output_7, label_9_input_7, 
      label_9_input_state_machine_7, nx5290, nx5294, nx5312, 
      label_9_output_8, label_9_input_8, label_9_input_state_machine_8, 
      nx18284, nx5322, nx5326, label_9_output_9, label_9_input_9, 
      label_9_input_state_machine_9, nx5354, nx5358, nx5376, 
      label_9_output_10, label_9_input_10, label_9_input_state_machine_10, 
      nx18287, nx5386, nx5390, label_9_output_11, label_9_input_11, 
      label_9_input_state_machine_11, nx5418, nx5422, nx5440, 
      label_9_output_12, label_9_input_12, label_9_input_state_machine_12, 
      nx18291, nx5450, nx5454, label_9_output_13, label_9_input_13, 
      label_9_input_state_machine_13, nx5482, nx5486, nx5504, nx5506, nx5508, 
      nx5512, nx5532, max_calc_comparator_fifth_inp2_13, 
      max_calc_comparator_fifth_inp1_13, max_calc_comparator_fifth_inp1_12, 
      nx5568, max_calc_comparator_fifth_inp2_11, 
      max_calc_comparator_fifth_inp1_11, max_calc_comparator_fifth_inp1_10, 
      nx5604, max_calc_comparator_fifth_inp2_9, 
      max_calc_comparator_fifth_inp1_9, max_calc_comparator_fifth_inp1_8, 
      nx5640, max_calc_comparator_fifth_inp2_7, 
      max_calc_comparator_fifth_inp1_7, max_calc_comparator_fifth_inp1_6, 
      nx5676, max_calc_comparator_fifth_inp2_5, 
      max_calc_comparator_fifth_inp1_5, max_calc_comparator_fifth_inp1_4, 
      nx5712, max_calc_comparator_fifth_inp2_3, 
      max_calc_comparator_fifth_inp1_3, max_calc_comparator_fifth_inp1_2, 
      nx5748, max_calc_comparator_fifth_inp2_1, nx5766, nx5790, nx5806, 
      nx5822, nx5838, nx5854, nx5870, nx5886, label_10_output_15, 
      label_10_input_15, label_10_input_state_machine_15, nx5910, nx5912, 
      nx5916, label_9_output_15, label_9_input_15, 
      label_9_input_state_machine_15, nx5950, nx5952, nx5956, nx5976, nx5978, 
      nx5986, nx5996, nx6000, max_calc_comparator_first_inp2_14, 
      label_2_output_14, label_2_input_14, label_2_input_state_machine_14, 
      label_2_output_0, label_2_input_0, booth_booth_integration_output_1_12, 
      booth_booth_integrtaion_1_shift_reg_output_9, 
      booth_booth_integrtaion_1_shift_Reg_count_9, output_8_dup_12716, 
      booth_booth_integrtaion_1_shift_Reg_count_8, output_7_dup_12717, 
      booth_booth_integrtaion_1_shift_Reg_count_7, output_6_dup_12718, 
      booth_booth_integrtaion_1_shift_Reg_count_6, output_5_dup_12719, 
      booth_booth_integrtaion_1_shift_Reg_count_5, output_4_dup_12720, 
      booth_booth_integrtaion_1_shift_Reg_count_4, output_3_dup_12721, 
      booth_booth_integrtaion_1_shift_Reg_count_3, output_2_dup_12722, 
      booth_booth_integrtaion_1_shift_Reg_count_2, output_1_dup_12723, 
      booth_booth_integrtaion_1_shift_Reg_count_1, 
      booth_booth_integrtaion_1_shift_reg_output_0, 
      booth_booth_integrtaion_1_shift_Reg_count_0, 
      booth_booth_integration_output_1_13, 
      booth_booth_integration_output_1_14, 
      booth_booth_integration_output_1_15, 
      booth_booth_integration_output_1_16, booth_output_0_dup_12130, 
      booth_output_1_dup_12129, booth_output_2_dup_12128, 
      booth_output_3_dup_12127, booth_output_4_dup_12126, 
      booth_output_5_dup_12125, booth_output_6_dup_12124, 
      booth_output_7_dup_12123, booth_output_8_dup_12122, 
      booth_output_9_dup_12121, booth_output_10_dup_12120, 
      booth_output_11_dup_12119, nx6108, nx6120, nx6132, nx6144, nx6156, 
      nx6168, nx6180, nx6192, nx6204, nx6216, nx6228, nx6240, nx6266, 
      booth_booth_integration_output_1_17, nx18297, nx6274, nx6280, nx6290, 
      booth_booth_integration_output_1_18, nx18299, nx6300, nx6304, nx6318, 
      booth_booth_integration_output_1_19, nx18300, nx6328, nx6338, 
      booth_booth_integration_output_1_20, nx18301, nx6348, nx6366, 
      booth_booth_integration_output_1_21, nx18302, nx6372, nx6376, nx6386, 
      booth_booth_integration_output_1_22, nx18303, nx6396, nx6414, 
      booth_booth_integration_output_1_23, nx18304, nx6420, nx6424, nx6434, 
      booth_booth_integration_output_1_24, nx18305, nx6444, nx6462, 
      booth_booth_integration_output_1_25, nx18307, nx6468, nx6472, nx6482, 
      booth_booth_integration_output_1_26, nx18309, nx6492, nx6510, 
      booth_booth_integration_output_1_27, nx18311, nx6516, nx6520, nx6530, 
      booth_output_28_dup_12118, nx18313, nx6540, nx6558, 
      booth_output_29_dup_12117, nx18315, nx6564, nx6568, nx6578, nx18317, 
      nx6588, nx6606, nx6614, nx6618, nx6630, nx6646, nx6654, nx6670, nx6678, 
      nx6694, nx6702, nx6718, nx6726, nx6742, nx6750, nx6762, nx6774, nx6790, 
      nx6796, nx6802, nx6820, nx6832, nx6844, nx6854, 
      label_2_input_state_machine_0, nx6866, label_2_output_1, 
      label_2_input_1, label_2_input_state_machine_1, nx6888, nx6892, nx6910, 
      label_2_output_2, label_2_input_2, label_2_input_state_machine_2, 
      nx18320, nx6920, nx6924, label_2_output_3, label_2_input_3, 
      label_2_input_state_machine_3, nx6952, nx6956, nx6974, 
      label_2_output_4, label_2_input_4, label_2_input_state_machine_4, 
      nx18322, nx6984, nx6988, label_2_output_5, label_2_input_5, 
      label_2_input_state_machine_5, nx7016, nx7020, nx7038, 
      label_2_output_6, label_2_input_6, label_2_input_state_machine_6, 
      nx18325, nx7048, nx7052, label_2_output_7, label_2_input_7, 
      label_2_input_state_machine_7, nx7080, nx7084, nx7102, 
      label_2_output_8, label_2_input_8, label_2_input_state_machine_8, 
      nx18329, nx7112, nx7116, label_2_output_9, label_2_input_9, 
      label_2_input_state_machine_9, nx7144, nx7148, nx7166, 
      label_2_output_10, label_2_input_10, label_2_input_state_machine_10, 
      nx18332, nx7176, nx7180, label_2_output_11, label_2_input_11, 
      label_2_input_state_machine_11, nx7208, nx7212, nx7230, 
      label_2_output_12, label_2_input_12, label_2_input_state_machine_12, 
      nx18334, nx7240, nx7244, label_2_output_13, label_2_input_13, 
      label_2_input_state_machine_13, nx7272, nx7276, nx7294, nx7296, nx7298, 
      nx7302, max_calc_ans2_14, max_calc_comparator_second_inp1_14, 
      label_3_output_14, label_3_input_14, label_3_input_state_machine_14, 
      label_3_output_0, label_3_input_0, booth_booth_integration_output_2_12, 
      booth_booth_integrtaion_2_shift_reg_output_9, 
      booth_booth_integrtaion_2_shift_Reg_count_9, output_8_dup_12744, 
      booth_booth_integrtaion_2_shift_Reg_count_8, output_7_dup_12745, 
      booth_booth_integrtaion_2_shift_Reg_count_7, output_6_dup_12746, 
      booth_booth_integrtaion_2_shift_Reg_count_6, output_5_dup_12747, 
      booth_booth_integrtaion_2_shift_Reg_count_5, output_4_dup_12748, 
      booth_booth_integrtaion_2_shift_Reg_count_4, output_3_dup_12749, 
      booth_booth_integrtaion_2_shift_Reg_count_3, output_2_dup_12750, 
      booth_booth_integrtaion_2_shift_Reg_count_2, output_1_dup_12751, 
      booth_booth_integrtaion_2_shift_Reg_count_1, 
      booth_booth_integrtaion_2_shift_reg_output_0, 
      booth_booth_integrtaion_2_shift_Reg_count_0, 
      booth_booth_integration_output_2_13, 
      booth_booth_integration_output_2_14, 
      booth_booth_integration_output_2_15, 
      booth_booth_integration_output_2_16, booth_output_0_dup_12149, 
      booth_output_1_dup_12148, booth_output_2_dup_12147, 
      booth_output_3_dup_12146, booth_output_4_dup_12145, 
      booth_output_5_dup_12144, booth_output_6_dup_12143, 
      booth_output_7_dup_12142, booth_output_8_dup_12141, 
      booth_output_9_dup_12140, booth_output_10_dup_12139, 
      booth_output_11_dup_12138, nx7418, nx7430, nx7442, nx7454, nx7466, 
      nx7478, nx7490, nx7502, nx7514, nx7526, nx7538, nx7550, nx7576, 
      booth_booth_integration_output_2_17, nx18337, nx7584, nx7590, nx7600, 
      booth_booth_integration_output_2_18, nx18339, nx7610, nx7614, nx7628, 
      booth_booth_integration_output_2_19, nx18341, nx7638, nx7648, 
      booth_booth_integration_output_2_20, nx18343, nx7658, nx7676, 
      booth_booth_integration_output_2_21, nx18345, nx7682, nx7686, nx7696, 
      booth_booth_integration_output_2_22, nx18347, nx7706, nx7724, 
      booth_booth_integration_output_2_23, nx18349, nx7730, nx7734, nx7744, 
      booth_booth_integration_output_2_24, nx18350, nx7754, nx7772, 
      booth_booth_integration_output_2_25, nx18351, nx7778, nx7782, nx7792, 
      booth_booth_integration_output_2_26, nx18352, nx7802, nx7820, 
      booth_booth_integration_output_2_27, nx18353, nx7826, nx7830, nx7840, 
      booth_output_28_dup_12137, nx18354, nx7850, nx7868, 
      booth_output_29_dup_12136, nx18355, nx7874, nx7878, nx7888, nx18357, 
      nx7898, nx7916, nx7924, nx7928, nx7940, nx7956, nx7964, nx7980, nx7988, 
      nx8004, nx8012, nx8028, nx8036, nx8052, nx8060, nx8072, nx8084, nx8100, 
      nx8106, nx8112, nx8130, nx8142, nx8154, nx8164, 
      label_3_input_state_machine_0, nx8176, label_3_output_1, 
      label_3_input_1, label_3_input_state_machine_1, nx8198, nx8202, nx8220, 
      label_3_output_2, label_3_input_2, label_3_input_state_machine_2, 
      nx18363, nx8230, nx8234, label_3_output_3, label_3_input_3, 
      label_3_input_state_machine_3, nx8262, nx8266, nx8284, 
      label_3_output_4, label_3_input_4, label_3_input_state_machine_4, 
      nx18365, nx8294, nx8298, label_3_output_5, label_3_input_5, 
      label_3_input_state_machine_5, nx8326, nx8330, nx8348, 
      label_3_output_6, label_3_input_6, label_3_input_state_machine_6, 
      nx18367, nx8358, nx8362, label_3_output_7, label_3_input_7, 
      label_3_input_state_machine_7, nx8390, nx8394, nx8412, 
      label_3_output_8, label_3_input_8, label_3_input_state_machine_8, 
      nx18369, nx8422, nx8426, label_3_output_9, label_3_input_9, 
      label_3_input_state_machine_9, nx8454, nx8458, nx8476, 
      label_3_output_10, label_3_input_10, label_3_input_state_machine_10, 
      nx18373, nx8486, nx8490, label_3_output_11, label_3_input_11, 
      label_3_input_state_machine_11, nx8518, nx8522, nx8540, 
      label_3_output_12, label_3_input_12, label_3_input_state_machine_12, 
      nx18376, nx8550, nx8554, label_3_output_13, label_3_input_13, 
      label_3_input_state_machine_13, nx8582, nx8586, nx8604, nx8606, nx8608, 
      nx8612, max_calc_ans3_14, max_calc_comparator_third_inp1_14, 
      label_5_output_14, label_5_input_14, label_5_input_state_machine_14, 
      label_5_output_0, label_5_input_0, booth_booth_integration_output_4_12, 
      booth_booth_integrtaion_4_shift_reg_output_9, 
      booth_booth_integrtaion_4_shift_Reg_count_9, output_8_dup_12800, 
      booth_booth_integrtaion_4_shift_Reg_count_8, output_7_dup_12801, 
      booth_booth_integrtaion_4_shift_Reg_count_7, output_6_dup_12802, 
      booth_booth_integrtaion_4_shift_Reg_count_6, output_5_dup_12803, 
      booth_booth_integrtaion_4_shift_Reg_count_5, output_4_dup_12804, 
      booth_booth_integrtaion_4_shift_Reg_count_4, output_3_dup_12805, 
      booth_booth_integrtaion_4_shift_Reg_count_3, output_2_dup_12806, 
      booth_booth_integrtaion_4_shift_Reg_count_2, output_1_dup_12807, 
      booth_booth_integrtaion_4_shift_Reg_count_1, 
      booth_booth_integrtaion_4_shift_reg_output_0, 
      booth_booth_integrtaion_4_shift_Reg_count_0, 
      booth_booth_integration_output_4_13, 
      booth_booth_integration_output_4_14, 
      booth_booth_integration_output_4_15, 
      booth_booth_integration_output_4_16, booth_output_0_dup_12187, 
      booth_output_1_dup_12186, booth_output_2_dup_12185, 
      booth_output_3_dup_12184, booth_output_4_dup_12183, 
      booth_output_5_dup_12182, booth_output_6_dup_12181, 
      booth_output_7_dup_12180, booth_output_8_dup_12179, 
      booth_output_9_dup_12178, booth_output_10_dup_12177, 
      booth_output_11_dup_12176, nx8738, nx8750, nx8762, nx8774, nx8786, 
      nx8798, nx8810, nx8822, nx8834, nx8846, nx8858, nx8870, nx8896, 
      booth_booth_integration_output_4_17, nx18379, nx8904, nx8910, nx8920, 
      booth_booth_integration_output_4_18, nx18380, nx8930, nx8934, nx8948, 
      booth_booth_integration_output_4_19, nx18381, nx8958, nx8968, 
      booth_booth_integration_output_4_20, nx18382, nx8978, nx8996, 
      booth_booth_integration_output_4_21, nx18383, nx9002, nx9006, nx9016, 
      booth_booth_integration_output_4_22, nx18385, nx9026, nx9044, 
      booth_booth_integration_output_4_23, nx18386, nx9050, nx9054, nx9064, 
      booth_booth_integration_output_4_24, nx18387, nx9074, nx9092, 
      booth_booth_integration_output_4_25, nx18388, nx9098, nx9102, nx9112, 
      booth_booth_integration_output_4_26, nx18389, nx9122, nx9140, 
      booth_booth_integration_output_4_27, nx18390, nx9146, nx9150, nx9160, 
      booth_output_28_dup_12175, nx18391, nx9170, nx9188, 
      booth_output_29_dup_12174, nx18393, nx9194, nx9198, nx9208, nx18395, 
      nx9218, nx9236, nx9244, nx9248, nx9260, nx9276, nx9284, nx9300, nx9308, 
      nx9324, nx9332, nx9348, nx9356, nx9372, nx9380, nx9392, nx9404, nx9420, 
      nx9426, nx9432, nx9450, nx9462, nx9474, nx9484, 
      label_5_input_state_machine_0, nx9496, label_5_output_1, 
      label_5_input_1, label_5_input_state_machine_1, nx9518, nx9522, nx9540, 
      label_5_output_2, label_5_input_2, label_5_input_state_machine_2, 
      nx18401, nx9550, nx9554, label_5_output_3, label_5_input_3, 
      label_5_input_state_machine_3, nx9582, nx9586, nx9604, 
      label_5_output_4, label_5_input_4, label_5_input_state_machine_4, 
      nx18403, nx9614, nx9618, label_5_output_5, label_5_input_5, 
      label_5_input_state_machine_5, nx9646, nx9650, nx9668, 
      label_5_output_6, label_5_input_6, label_5_input_state_machine_6, 
      nx18405, nx9678, nx9682, label_5_output_7, label_5_input_7, 
      label_5_input_state_machine_7, nx9710, nx9714, nx9732, 
      label_5_output_8, label_5_input_8, label_5_input_state_machine_8, 
      nx18407, nx9742, nx9746, label_5_output_9, label_5_input_9, 
      label_5_input_state_machine_9, nx9774, nx9778, nx9796, 
      label_5_output_10, label_5_input_10, label_5_input_state_machine_10, 
      nx18411, nx9806, nx9810, label_5_output_11, label_5_input_11, 
      label_5_input_state_machine_11, nx9838, nx9842, nx9860, 
      label_5_output_12, label_5_input_12, label_5_input_state_machine_12, 
      nx18415, nx9870, nx9874, label_5_output_13, label_5_input_13, 
      label_5_input_state_machine_13, nx9902, nx9906, nx9924, nx9926, nx9928, 
      nx9932, label_6_output_14, label_6_input_14, 
      label_6_input_state_machine_14, label_6_output_0, label_6_input_0, 
      booth_booth_integration_output_5_12, 
      booth_booth_integrtaion_5_shift_reg_output_9, 
      booth_booth_integrtaion_5_shift_Reg_count_9, output_8_dup_12828, 
      booth_booth_integrtaion_5_shift_Reg_count_8, output_7_dup_12829, 
      booth_booth_integrtaion_5_shift_Reg_count_7, output_6_dup_12830, 
      booth_booth_integrtaion_5_shift_Reg_count_6, output_5_dup_12831, 
      booth_booth_integrtaion_5_shift_Reg_count_5, output_4_dup_12832, 
      booth_booth_integrtaion_5_shift_Reg_count_4, output_3_dup_12833, 
      booth_booth_integrtaion_5_shift_Reg_count_3, output_2_dup_12834, 
      booth_booth_integrtaion_5_shift_Reg_count_2, output_1_dup_12835, 
      booth_booth_integrtaion_5_shift_Reg_count_1, 
      booth_booth_integrtaion_5_shift_reg_output_0, 
      booth_booth_integrtaion_5_shift_Reg_count_0, 
      booth_booth_integration_output_5_13, 
      booth_booth_integration_output_5_14, 
      booth_booth_integration_output_5_15, 
      booth_booth_integration_output_5_16, booth_output_0_dup_12206, 
      booth_output_1_dup_12205, booth_output_2_dup_12204, 
      booth_output_3_dup_12203, booth_output_4_dup_12202, 
      booth_output_5_dup_12201, booth_output_6_dup_12200, 
      booth_output_7_dup_12199, booth_output_8_dup_12198, 
      booth_output_9_dup_12197, booth_output_10_dup_12196, 
      booth_output_11_dup_12195, nx10056, nx10068, nx10080, nx10092, nx10104, 
      nx10116, nx10128, nx10140, nx10152, nx10164, nx10176, nx10188, nx10214, 
      booth_booth_integration_output_5_17, nx18421, nx10222, nx10228, 
      nx10238, booth_booth_integration_output_5_18, nx18422, nx10248, 
      nx10252, nx10266, booth_booth_integration_output_5_19, nx18423, 
      nx10276, nx10286, booth_booth_integration_output_5_20, nx18424, 
      nx10296, nx10314, booth_booth_integration_output_5_21, nx18425, 
      nx10320, nx10324, nx10334, booth_booth_integration_output_5_22, 
      nx18426, nx10344, nx10362, booth_booth_integration_output_5_23, 
      nx18427, nx10368, nx10372, nx10382, 
      booth_booth_integration_output_5_24, nx18429, nx10392, nx10410, 
      booth_booth_integration_output_5_25, nx18431, nx10416, nx10420, 
      nx10430, booth_booth_integration_output_5_26, nx18433, nx10440, 
      nx10458, booth_booth_integration_output_5_27, nx18435, nx10464, 
      nx10468, nx10478, booth_output_28_dup_12194, nx18437, nx10488, nx10506, 
      booth_output_29_dup_12193, nx18439, nx10512, nx10516, nx10526, nx18440, 
      nx10536, nx10554, nx10562, nx10566, nx10578, nx10594, nx10602, nx10618, 
      nx10626, nx10642, nx10650, nx10666, nx10674, nx10690, nx10698, nx10710, 
      nx10722, nx10738, nx10744, nx10750, nx10768, nx10780, nx10792, nx10802, 
      label_6_input_state_machine_0, nx10814, label_6_output_1, 
      label_6_input_1, label_6_input_state_machine_1, nx10836, nx10840, 
      nx10858, label_6_output_2, label_6_input_2, 
      label_6_input_state_machine_2, nx18443, nx10868, nx10872, 
      label_6_output_3, label_6_input_3, label_6_input_state_machine_3, 
      nx10900, nx10904, nx10922, label_6_output_4, label_6_input_4, 
      label_6_input_state_machine_4, nx18445, nx10932, nx10936, 
      label_6_output_5, label_6_input_5, label_6_input_state_machine_5, 
      nx10964, nx10968, nx10986, label_6_output_6, label_6_input_6, 
      label_6_input_state_machine_6, nx18449, nx10996, nx11000, 
      label_6_output_7, label_6_input_7, label_6_input_state_machine_7, 
      nx11028, nx11032, nx11050, label_6_output_8, label_6_input_8, 
      label_6_input_state_machine_8, nx18453, nx11060, nx11064, 
      label_6_output_9, label_6_input_9, label_6_input_state_machine_9, 
      nx11092, nx11096, nx11114, label_6_output_10, label_6_input_10, 
      label_6_input_state_machine_10, nx18455, nx11124, nx11128, 
      label_6_output_11, label_6_input_11, label_6_input_state_machine_11, 
      nx11156, nx11160, nx11178, label_6_output_12, label_6_input_12, 
      label_6_input_state_machine_12, nx18457, nx11188, nx11192, 
      label_6_output_13, label_6_input_13, label_6_input_state_machine_13, 
      nx11220, nx11224, nx11242, nx11244, nx11246, nx11250, nx11272, 
      max_calc_comparator_third_inp2_13, max_calc_comparator_third_inp1_13, 
      max_calc_comparator_third_inp1_12, nx11316, 
      max_calc_comparator_third_inp2_11, max_calc_comparator_third_inp1_11, 
      max_calc_comparator_third_inp1_10, nx11360, 
      max_calc_comparator_third_inp2_9, max_calc_comparator_third_inp1_9, 
      max_calc_comparator_third_inp1_8, nx11404, 
      max_calc_comparator_third_inp2_7, max_calc_comparator_third_inp1_7, 
      max_calc_comparator_third_inp1_6, nx11448, 
      max_calc_comparator_third_inp2_5, max_calc_comparator_third_inp1_5, 
      max_calc_comparator_third_inp1_4, nx11492, 
      max_calc_comparator_third_inp2_3, max_calc_comparator_third_inp1_3, 
      max_calc_comparator_third_inp1_2, nx11536, 
      max_calc_comparator_third_inp2_1, nx11558, 
      max_calc_comparator_third_inp1_0, nx11594, nx11610, nx11626, nx11642, 
      nx11658, nx11674, nx11690, label_6_output_15, label_6_input_15, 
      label_6_input_state_machine_15, nx11714, nx11716, nx11720, 
      label_5_output_15, label_5_input_15, label_5_input_state_machine_15, 
      nx11756, nx11758, nx11762, nx11784, nx11786, nx11794, nx11808, 
      label_4_output_14, label_4_input_14, label_4_input_state_machine_14, 
      label_4_output_0, label_4_input_0, booth_booth_integration_output_3_12, 
      booth_booth_integrtaion_3_shift_reg_output_9, 
      booth_booth_integrtaion_3_shift_Reg_count_9, output_8_dup_12772, 
      booth_booth_integrtaion_3_shift_Reg_count_8, output_7_dup_12773, 
      booth_booth_integrtaion_3_shift_Reg_count_7, output_6_dup_12774, 
      booth_booth_integrtaion_3_shift_Reg_count_6, output_5_dup_12775, 
      booth_booth_integrtaion_3_shift_Reg_count_5, output_4_dup_12776, 
      booth_booth_integrtaion_3_shift_Reg_count_4, output_3_dup_12777, 
      booth_booth_integrtaion_3_shift_Reg_count_3, output_2_dup_12778, 
      booth_booth_integrtaion_3_shift_Reg_count_2, output_1_dup_12779, 
      booth_booth_integrtaion_3_shift_Reg_count_1, 
      booth_booth_integrtaion_3_shift_reg_output_0, 
      booth_booth_integrtaion_3_shift_Reg_count_0, 
      booth_booth_integration_output_3_13, 
      booth_booth_integration_output_3_14, 
      booth_booth_integration_output_3_15, 
      booth_booth_integration_output_3_16, booth_output_0_dup_12168, 
      booth_output_1_dup_12167, booth_output_2_dup_12166, 
      booth_output_3_dup_12165, booth_output_4_dup_12164, 
      booth_output_5_dup_12163, booth_output_6_dup_12162, 
      booth_output_7_dup_12161, booth_output_8_dup_12160, 
      booth_output_9_dup_12159, booth_output_10_dup_12158, 
      booth_output_11_dup_12157, nx11920, nx11932, nx11944, nx11956, nx11968, 
      nx11980, nx11992, nx12004, nx12016, nx12028, nx12040, nx12052, nx12078, 
      booth_booth_integration_output_3_17, nx18461, nx12086, nx12092, 
      nx12102, booth_booth_integration_output_3_18, nx18463, nx12112, 
      nx12116, nx12130, booth_booth_integration_output_3_19, nx18465, 
      nx12140, nx12150, booth_booth_integration_output_3_20, nx18467, 
      nx12160, nx12178, booth_booth_integration_output_3_21, nx18469, 
      nx12184, nx12188, nx12198, booth_booth_integration_output_3_22, 
      nx18471, nx12208, nx12226, booth_booth_integration_output_3_23, 
      nx18472, nx12232, nx12236, nx12246, 
      booth_booth_integration_output_3_24, nx18473, nx12256, nx12274, 
      booth_booth_integration_output_3_25, nx18474, nx12280, nx12284, 
      nx12294, booth_booth_integration_output_3_26, nx18475, nx12304, 
      nx12322, booth_booth_integration_output_3_27, nx18476, nx12328, 
      nx12332, nx12342, booth_output_28_dup_12156, nx18477, nx12352, nx12370, 
      booth_output_29_dup_12155, nx18479, nx12376, nx12380, nx12390, nx18481, 
      nx12400, nx12418, nx12426, nx12430, nx12442, nx12458, nx12466, nx12482, 
      nx12490, nx12506, nx12514, nx12530, nx12538, nx12554, nx12562, nx12574, 
      nx12586, nx12602, nx12608, nx12614, nx12632, nx12644, nx12656, nx12666, 
      label_4_input_state_machine_0, nx12678, label_4_output_1, 
      label_4_input_1, label_4_input_state_machine_1, nx12700, nx12704, 
      nx12722, label_4_output_2, label_4_input_2, 
      label_4_input_state_machine_2, nx18486, nx12732, nx12736, 
      label_4_output_3, label_4_input_3, label_4_input_state_machine_3, 
      nx12764, nx12768, nx12786, label_4_output_4, label_4_input_4, 
      label_4_input_state_machine_4, nx18488, nx12796, nx12800, 
      label_4_output_5, label_4_input_5, label_4_input_state_machine_5, 
      nx12828, nx12832, nx12850, label_4_output_6, label_4_input_6, 
      label_4_input_state_machine_6, nx18490, nx12860, nx12864, 
      label_4_output_7, label_4_input_7, label_4_input_state_machine_7, 
      nx12892, nx12896, nx12914, label_4_output_8, label_4_input_8, 
      label_4_input_state_machine_8, nx18493, nx12924, nx12928, 
      label_4_output_9, label_4_input_9, label_4_input_state_machine_9, 
      nx12956, nx12960, nx12978, label_4_output_10, label_4_input_10, 
      label_4_input_state_machine_10, nx18497, nx12988, nx12992, 
      label_4_output_11, label_4_input_11, label_4_input_state_machine_11, 
      nx13020, nx13024, nx13042, label_4_output_12, label_4_input_12, 
      label_4_input_state_machine_12, nx18499, nx13052, nx13056, 
      label_4_output_13, label_4_input_13, label_4_input_state_machine_13, 
      nx13084, nx13088, nx13106, nx13108, nx13110, nx13114, max_calc_ans4_14, 
      max_calc_comparator_fourth_inp1_14, label_7_output_14, 
      label_7_input_14, label_7_input_state_machine_14, label_7_output_0, 
      label_7_input_0, booth_booth_integration_output_6_12, 
      booth_booth_integrtaion_6_shift_reg_output_9, 
      booth_booth_integrtaion_6_shift_Reg_count_9, output_8_dup_12856, 
      booth_booth_integrtaion_6_shift_Reg_count_8, output_7_dup_12857, 
      booth_booth_integrtaion_6_shift_Reg_count_7, output_6_dup_12858, 
      booth_booth_integrtaion_6_shift_Reg_count_6, output_5_dup_12859, 
      booth_booth_integrtaion_6_shift_Reg_count_5, output_4_dup_12860, 
      booth_booth_integrtaion_6_shift_Reg_count_4, output_3_dup_12861, 
      booth_booth_integrtaion_6_shift_Reg_count_3, output_2_dup_12862, 
      booth_booth_integrtaion_6_shift_Reg_count_2, output_1_dup_12863, 
      booth_booth_integrtaion_6_shift_Reg_count_1, 
      booth_booth_integrtaion_6_shift_reg_output_0, 
      booth_booth_integrtaion_6_shift_Reg_count_0, 
      booth_booth_integration_output_6_13, 
      booth_booth_integration_output_6_14, 
      booth_booth_integration_output_6_15, 
      booth_booth_integration_output_6_16, booth_output_0_dup_12225, 
      booth_output_1_dup_12224, booth_output_2_dup_12223, 
      booth_output_3_dup_12222, booth_output_4_dup_12221, 
      booth_output_5_dup_12220, booth_output_6_dup_12219, 
      booth_output_7_dup_12218, booth_output_8_dup_12217, 
      booth_output_9_dup_12216, booth_output_10_dup_12215, 
      booth_output_11_dup_12214, nx13230, nx13242, nx13254, nx13266, nx13278, 
      nx13290, nx13302, nx13314, nx13326, nx13338, nx13350, nx13362, nx13388, 
      booth_booth_integration_output_6_17, nx18502, nx13396, nx13402, 
      nx13412, booth_booth_integration_output_6_18, nx18503, nx13422, 
      nx13426, nx13440, booth_booth_integration_output_6_19, nx18504, 
      nx13450, nx13460, booth_booth_integration_output_6_20, nx18505, 
      nx13470, nx13488, booth_booth_integration_output_6_21, nx18507, 
      nx13494, nx13498, nx13508, booth_booth_integration_output_6_22, 
      nx18508, nx13518, nx13536, booth_booth_integration_output_6_23, 
      nx18509, nx13542, nx13546, nx13556, 
      booth_booth_integration_output_6_24, nx18510, nx13566, nx13584, 
      booth_booth_integration_output_6_25, nx18511, nx13590, nx13594, 
      nx13604, booth_booth_integration_output_6_26, nx18512, nx13614, 
      nx13632, booth_booth_integration_output_6_27, nx18513, nx13638, 
      nx13642, nx13652, booth_output_28_dup_12213, nx18515, nx13662, nx13680, 
      booth_output_29_dup_12212, nx18517, nx13686, nx13690, nx13700, nx18519, 
      nx13710, nx13728, nx13736, nx13740, nx13752, nx13768, nx13776, nx13792, 
      nx13800, nx13816, nx13824, nx13840, nx13848, nx13864, nx13872, nx13884, 
      nx13896, nx13912, nx13918, nx13924, nx13942, nx13954, nx13966, nx13976, 
      label_7_input_state_machine_0, nx13988, label_7_output_1, 
      label_7_input_1, label_7_input_state_machine_1, nx14010, nx14014, 
      nx14032, label_7_output_2, label_7_input_2, 
      label_7_input_state_machine_2, nx18524, nx14042, nx14046, 
      label_7_output_3, label_7_input_3, label_7_input_state_machine_3, 
      nx14074, nx14078, nx14096, label_7_output_4, label_7_input_4, 
      label_7_input_state_machine_4, nx18526, nx14106, nx14110, 
      label_7_output_5, label_7_input_5, label_7_input_state_machine_5, 
      nx14138, nx14142, nx14160, label_7_output_6, label_7_input_6, 
      label_7_input_state_machine_6, nx18528, nx14170, nx14174, 
      label_7_output_7, label_7_input_7, label_7_input_state_machine_7, 
      nx14202, nx14206, nx14224, label_7_output_8, label_7_input_8, 
      label_7_input_state_machine_8, nx18531, nx14234, nx14238, 
      label_7_output_9, label_7_input_9, label_7_input_state_machine_9, 
      nx14266, nx14270, nx14288, label_7_output_10, label_7_input_10, 
      label_7_input_state_machine_10, nx18535, nx14298, nx14302, 
      label_7_output_11, label_7_input_11, label_7_input_state_machine_11, 
      nx14330, nx14334, nx14352, label_7_output_12, label_7_input_12, 
      label_7_input_state_machine_12, nx18539, nx14362, nx14366, 
      label_7_output_13, label_7_input_13, label_7_input_state_machine_13, 
      nx14394, nx14398, nx14416, nx14418, nx14420, nx14424, 
      label_8_output_14, label_8_input_14, label_8_input_state_machine_14, 
      label_8_output_0, label_8_input_0, booth_booth_integration_output_7_12, 
      booth_booth_integrtaion_7_shift_reg_output_9, 
      booth_booth_integrtaion_7_shift_Reg_count_9, output_8_dup_12884, 
      booth_booth_integrtaion_7_shift_Reg_count_8, output_7_dup_12885, 
      booth_booth_integrtaion_7_shift_Reg_count_7, output_6_dup_12886, 
      booth_booth_integrtaion_7_shift_Reg_count_6, output_5_dup_12887, 
      booth_booth_integrtaion_7_shift_Reg_count_5, output_4_dup_12888, 
      booth_booth_integrtaion_7_shift_Reg_count_4, output_3_dup_12889, 
      booth_booth_integrtaion_7_shift_Reg_count_3, output_2_dup_12890, 
      booth_booth_integrtaion_7_shift_Reg_count_2, output_1_dup_12891, 
      booth_booth_integrtaion_7_shift_Reg_count_1, 
      booth_booth_integrtaion_7_shift_reg_output_0, 
      booth_booth_integrtaion_7_shift_Reg_count_0, 
      booth_booth_integration_output_7_13, 
      booth_booth_integration_output_7_14, 
      booth_booth_integration_output_7_15, 
      booth_booth_integration_output_7_16, booth_output_0_dup_12244, 
      booth_output_1_dup_12243, booth_output_2_dup_12242, 
      booth_output_3_dup_12241, booth_output_4_dup_12240, 
      booth_output_5_dup_12239, booth_output_6_dup_12238, 
      booth_output_7_dup_12237, booth_output_8_dup_12236, 
      booth_output_9_dup_12235, booth_output_10_dup_12234, 
      booth_output_11_dup_12233, nx14546, nx14558, nx14570, nx14582, nx14594, 
      nx14606, nx14618, nx14630, nx14642, nx14654, nx14666, nx14678, nx14704, 
      booth_booth_integration_output_7_17, nx18544, nx14712, nx14718, 
      nx14728, booth_booth_integration_output_7_18, nx18545, nx14738, 
      nx14742, nx14756, booth_booth_integration_output_7_19, nx18546, 
      nx14766, nx14776, booth_booth_integration_output_7_20, nx18547, 
      nx14786, nx14804, booth_booth_integration_output_7_21, nx18548, 
      nx14810, nx14814, nx14824, booth_booth_integration_output_7_22, 
      nx18549, nx14834, nx14852, booth_booth_integration_output_7_23, 
      nx18551, nx14858, nx14862, nx14872, 
      booth_booth_integration_output_7_24, nx18553, nx14882, nx14900, 
      booth_booth_integration_output_7_25, nx18555, nx14906, nx14910, 
      nx14920, booth_booth_integration_output_7_26, nx18557, nx14930, 
      nx14948, booth_booth_integration_output_7_27, nx18559, nx14954, 
      nx14958, nx14968, booth_output_28_dup_12232, nx18561, nx14978, nx14996, 
      booth_output_29_dup_12231, nx18562, nx15002, nx15006, nx15016, nx18563, 
      nx15026, nx15044, nx15052, nx15056, nx15068, nx15084, nx15092, nx15108, 
      nx15116, nx15132, nx15140, nx15156, nx15164, nx15180, nx15188, nx15200, 
      nx15212, nx15228, nx15234, nx15240, nx15258, nx15270, nx15282, nx15292, 
      label_8_input_state_machine_0, nx15304, label_8_output_1, 
      label_8_input_1, label_8_input_state_machine_1, nx15326, nx15330, 
      nx15348, label_8_output_2, label_8_input_2, 
      label_8_input_state_machine_2, nx18566, nx15358, nx15362, 
      label_8_output_3, label_8_input_3, label_8_input_state_machine_3, 
      nx15390, nx15394, nx15412, label_8_output_4, label_8_input_4, 
      label_8_input_state_machine_4, nx18569, nx15422, nx15426, 
      label_8_output_5, label_8_input_5, label_8_input_state_machine_5, 
      nx15454, nx15458, nx15476, label_8_output_6, label_8_input_6, 
      label_8_input_state_machine_6, nx18573, nx15486, nx15490, 
      label_8_output_7, label_8_input_7, label_8_input_state_machine_7, 
      nx15518, nx15522, nx15540, label_8_output_8, label_8_input_8, 
      label_8_input_state_machine_8, nx18576, nx15550, nx15554, 
      label_8_output_9, label_8_input_9, label_8_input_state_machine_9, 
      nx15582, nx15586, nx15604, label_8_output_10, label_8_input_10, 
      label_8_input_state_machine_10, nx18578, nx15614, nx15618, 
      label_8_output_11, label_8_input_11, label_8_input_state_machine_11, 
      nx15646, nx15650, nx15668, label_8_output_12, label_8_input_12, 
      label_8_input_state_machine_12, nx18580, nx15678, nx15682, 
      label_8_output_13, label_8_input_13, label_8_input_state_machine_13, 
      nx15710, nx15714, nx15732, nx15734, nx15736, nx15740, nx15762, 
      max_calc_comparator_fourth_inp2_13, max_calc_comparator_fourth_inp1_13, 
      max_calc_comparator_fourth_inp1_12, nx15806, 
      max_calc_comparator_fourth_inp2_11, max_calc_comparator_fourth_inp1_11, 
      max_calc_comparator_fourth_inp1_10, nx15850, 
      max_calc_comparator_fourth_inp2_9, max_calc_comparator_fourth_inp1_9, 
      max_calc_comparator_fourth_inp1_8, nx15894, 
      max_calc_comparator_fourth_inp2_7, max_calc_comparator_fourth_inp1_7, 
      max_calc_comparator_fourth_inp1_6, nx15938, 
      max_calc_comparator_fourth_inp2_5, max_calc_comparator_fourth_inp1_5, 
      max_calc_comparator_fourth_inp1_4, nx15982, 
      max_calc_comparator_fourth_inp2_3, max_calc_comparator_fourth_inp1_3, 
      max_calc_comparator_fourth_inp1_2, nx16026, 
      max_calc_comparator_fourth_inp2_1, nx16048, 
      max_calc_comparator_fourth_inp1_0, nx16084, nx16100, nx16116, nx16132, 
      nx16148, nx16164, nx16180, label_8_output_15, label_8_input_15, 
      label_8_input_state_machine_15, nx16204, nx16206, nx16210, 
      label_7_output_15, label_7_input_15, label_7_input_state_machine_15, 
      nx16246, nx16248, nx16252, nx16274, nx16276, nx16284, nx16298, nx16310, 
      max_calc_comparator_second_inp2_13, max_calc_ans4_13, nx16322, nx16336, 
      max_calc_comparator_second_inp1_13, max_calc_ans3_13, nx16358, nx16372, 
      max_calc_ans4_12, nx16396, nx16410, max_calc_comparator_second_inp1_12, 
      max_calc_ans3_12, nx16432, nx16446, nx16458, 
      max_calc_comparator_second_inp2_11, max_calc_ans4_11, nx16470, nx16484, 
      max_calc_comparator_second_inp1_11, max_calc_ans3_11, nx16506, nx16520, 
      max_calc_ans4_10, nx16544, nx16558, max_calc_comparator_second_inp1_10, 
      max_calc_ans3_10, nx16580, nx16594, nx16606, 
      max_calc_comparator_second_inp2_9, max_calc_ans4_9, nx16618, nx16632, 
      max_calc_comparator_second_inp1_9, max_calc_ans3_9, nx16654, nx16668, 
      max_calc_ans4_8, nx16692, nx16706, max_calc_comparator_second_inp1_8, 
      max_calc_ans3_8, nx16728, nx16742, nx16754, 
      max_calc_comparator_second_inp2_7, max_calc_ans4_7, nx16766, nx16780, 
      max_calc_comparator_second_inp1_7, max_calc_ans3_7, nx16802, nx16816, 
      max_calc_ans4_6, nx16840, nx16854, max_calc_comparator_second_inp1_6, 
      max_calc_ans3_6, nx16876, nx16890, nx16902, 
      max_calc_comparator_second_inp2_5, max_calc_ans4_5, nx16914, nx16928, 
      max_calc_comparator_second_inp1_5, max_calc_ans3_5, nx16950, nx16964, 
      max_calc_ans4_4, nx16988, nx17002, max_calc_comparator_second_inp1_4, 
      max_calc_ans3_4, nx17024, nx17038, nx17050, 
      max_calc_comparator_second_inp2_3, max_calc_ans4_3, nx17062, nx17076, 
      max_calc_comparator_second_inp1_3, max_calc_ans3_3, nx17098, nx17112, 
      max_calc_ans4_2, nx17136, nx17150, max_calc_comparator_second_inp1_2, 
      max_calc_ans3_2, nx17172, nx17186, nx17198, 
      max_calc_comparator_second_inp2_1, max_calc_ans4_1, nx17210, nx17224, 
      max_calc_ans3_1, nx17246, nx17260, nx17272, max_calc_ans4_0, nx17284, 
      nx17298, max_calc_comparator_second_inp1_0, max_calc_ans3_0, nx17320, 
      nx17334, nx17360, nx17376, nx17392, nx17408, nx17424, nx17440, nx17456, 
      label_4_output_15, label_4_input_15, label_4_input_state_machine_15, 
      nx17480, nx17482, nx17486, max_calc_ans4_15, nx17508, nx17522, 
      label_3_output_15, label_3_input_15, label_3_input_state_machine_15, 
      nx17548, nx17550, nx17554, max_calc_ans3_15, nx17576, nx17590, nx17602, 
      nx17604, nx17612, nx17622, max_calc_ans8_14, 
      max_calc_comparator_first_inp1_14, label_1_output_14, label_1_input_14, 
      label_1_input_state_machine_14, label_1_output_1, label_1_input_1, 
      label_1_input_state_machine_1, nx17644, nx17648, nx17666, 
      label_1_output_2, label_1_input_2, label_1_input_state_machine_2, 
      nx18585, nx17676, nx17680, label_1_output_3, label_1_input_3, 
      label_1_input_state_machine_3, nx17708, nx17712, nx17730, 
      label_1_output_4, label_1_input_4, label_1_input_state_machine_4, 
      nx18589, nx17740, nx17744, label_1_output_5, label_1_input_5, 
      label_1_input_state_machine_5, nx17772, nx17776, nx17794, 
      label_1_output_6, label_1_input_6, label_1_input_state_machine_6, 
      nx18593, nx17804, nx17808, label_1_output_7, label_1_input_7, 
      label_1_input_state_machine_7, nx17836, nx17840, nx17858, 
      label_1_output_8, label_1_input_8, label_1_input_state_machine_8, 
      nx18595, nx17868, nx17872, label_1_output_9, label_1_input_9, 
      label_1_input_state_machine_9, nx17900, nx17904, nx17922, 
      label_1_output_10, label_1_input_10, label_1_input_state_machine_10, 
      nx18597, nx17932, nx17936, label_1_output_11, label_1_input_11, 
      label_1_input_state_machine_11, nx17964, nx17968, nx17986, 
      label_1_output_12, label_1_input_12, label_1_input_state_machine_12, 
      nx18599, nx17996, nx18000, label_1_output_13, label_1_input_13, 
      label_1_input_state_machine_13, nx18028, nx18032, nx18050, nx18052, 
      nx18054, nx18058, max_calc_ans1_14, nx18603, nx18082, max_calc_ans6_14, 
      max_calc_ans5_14, nx18104, nx18114, nx18118, nx18605, max_calc_ans7_14, 
      nx18152, nx18156, nx18164, max_calc_comparator_first_inp2_13, 
      max_calc_ans2_13, nx18176, nx18186, max_calc_ans8_13, 
      max_calc_comparator_first_inp1_13, max_calc_ans1_13, nx18607, nx18204, 
      max_calc_ans6_13, max_calc_ans5_13, nx18226, nx18236, nx18240, 
      max_calc_ans7_13, nx18274, nx18278, max_calc_comparator_first_inp2_12, 
      max_calc_ans2_12, nx18298, nx18308, max_calc_ans8_12, 
      max_calc_comparator_first_inp1_12, max_calc_ans1_12, nx18608, nx18326, 
      max_calc_ans6_12, max_calc_ans5_12, nx18348, nx18358, nx18362, 
      max_calc_ans7_12, nx18396, nx18400, nx18408, 
      max_calc_comparator_first_inp2_11, max_calc_ans2_11, nx18420, nx18430, 
      max_calc_ans8_11, max_calc_comparator_first_inp1_11, max_calc_ans1_11, 
      nx18609, nx18448, max_calc_ans6_11, max_calc_ans5_11, nx18470, nx18480, 
      nx18484, max_calc_ans7_11, nx18518, nx18522, 
      max_calc_comparator_first_inp2_10, max_calc_ans2_10, nx18542, nx18552, 
      max_calc_ans8_10, max_calc_comparator_first_inp1_10, max_calc_ans1_10, 
      nx18610, nx18570, max_calc_ans6_10, max_calc_ans5_10, nx18592, nx18602, 
      nx18606, max_calc_ans7_10, nx18640, nx18644, nx18652, 
      max_calc_comparator_first_inp2_9, max_calc_ans2_9, nx18664, nx18674, 
      max_calc_ans8_9, max_calc_comparator_first_inp1_9, max_calc_ans1_9, 
      nx18611, nx18692, max_calc_ans6_9, max_calc_ans5_9, nx18714, nx18724, 
      nx18728, max_calc_ans7_9, nx18762, nx18766, 
      max_calc_comparator_first_inp2_8, max_calc_ans2_8, nx18786, nx18796, 
      max_calc_ans8_8, max_calc_comparator_first_inp1_8, max_calc_ans1_8, 
      nx18612, nx18814, max_calc_ans6_8, max_calc_ans5_8, nx18836, nx18846, 
      nx18850, max_calc_ans7_8, nx18884, nx18888, nx18896, 
      max_calc_comparator_first_inp2_7, max_calc_ans2_7, nx18908, nx18918, 
      max_calc_ans8_7, max_calc_comparator_first_inp1_7, max_calc_ans1_7, 
      nx18613, nx18936, max_calc_ans6_7, max_calc_ans5_7, nx18958, nx18968, 
      nx18972, max_calc_ans7_7, nx19006, nx19010, 
      max_calc_comparator_first_inp2_6, max_calc_ans2_6, nx19030, nx19040, 
      max_calc_ans8_6, max_calc_comparator_first_inp1_6, max_calc_ans1_6, 
      nx18615, nx19058, max_calc_ans6_6, max_calc_ans5_6, nx19080, nx19090, 
      nx19094, max_calc_ans7_6, nx19128, nx19132, nx19140, 
      max_calc_comparator_first_inp2_5, max_calc_ans2_5, nx19152, nx19162, 
      max_calc_ans8_5, max_calc_comparator_first_inp1_5, max_calc_ans1_5, 
      nx18617, nx19180, max_calc_ans6_5, max_calc_ans5_5, nx19202, nx19212, 
      nx19216, max_calc_ans7_5, nx19250, nx19254, 
      max_calc_comparator_first_inp2_4, max_calc_ans2_4, nx19274, nx19284, 
      max_calc_ans8_4, max_calc_comparator_first_inp1_4, max_calc_ans1_4, 
      nx18619, nx19302, max_calc_ans6_4, max_calc_ans5_4, nx19324, nx19334, 
      nx19338, max_calc_ans7_4, nx19372, nx19376, nx19384, 
      max_calc_comparator_first_inp2_3, max_calc_ans2_3, nx19396, nx19406, 
      max_calc_ans8_3, max_calc_comparator_first_inp1_3, max_calc_ans1_3, 
      nx18620, nx19424, max_calc_ans6_3, max_calc_ans5_3, nx19446, nx19456, 
      nx19460, max_calc_ans7_3, nx19494, nx19498, 
      max_calc_comparator_first_inp2_2, max_calc_ans2_2, nx19518, nx19528, 
      max_calc_ans8_2, max_calc_comparator_first_inp1_2, max_calc_ans1_2, 
      nx18621, nx19546, max_calc_ans6_2, max_calc_ans5_2, nx19568, nx19578, 
      nx19582, max_calc_ans7_2, nx19616, nx19620, nx19628, 
      max_calc_comparator_first_inp2_1, max_calc_ans2_1, nx19640, nx19650, 
      max_calc_ans8_1, max_calc_comparator_first_inp1_1, max_calc_ans1_1, 
      nx18622, nx19668, max_calc_ans6_1, max_calc_ans5_1, nx19690, nx19700, 
      nx19704, max_calc_ans7_1, nx19738, nx19742, nx19750, 
      max_calc_comparator_first_inp2_0, max_calc_ans2_0, nx19762, nx19772, 
      max_calc_ans8_0, max_calc_ans7_0, nx19796, nx19800, nx19822, nx19838, 
      nx19854, nx19870, nx19886, nx19902, nx19918, 
      max_calc_comparator_first_inp2_15, label_2_output_15, label_2_input_15, 
      label_2_input_state_machine_15, nx19942, nx19944, nx19948, 
      max_calc_ans2_15, nx19970, nx19980, max_calc_ans8_15, 
      max_calc_comparator_first_inp1_15, label_1_output_15, label_1_input_15, 
      label_1_input_state_machine_15, nx20000, nx20002, nx20006, 
      max_calc_ans1_15, nx18623, nx20030, max_calc_ans6_15, max_calc_ans5_15, 
      nx20052, nx20062, nx20066, max_calc_ans7_15, nx20100, nx20104, nx20112, 
      max_calc_answer_1, max_calc_answer_2, max_calc_answer_3, nx20152, 
      max_calc_answer_4, max_calc_answer_5, max_calc_answer_6, 
      max_calc_answer_7, nx20182, max_calc_answer_8, max_calc_answer_9, 
      max_calc_answer_10, max_calc_answer_11, nx20214, max_calc_answer_12, 
      max_calc_answer_13, max_calc_answer_14, max_calc_answer_15, nx20244, 
      nx20262, nx20276, nx20292, nx20306, nx20324, nx20338, nx20354, nx20368, 
      nx20386, nx20400, nx20416, nx20430, nx20448, nx20462, nx20478, nx20492, 
      nx20510, nx20524, nx20540, nx20554, nx20558, nx20652, nx20664, nx20758, 
      nx20772, nx20786, nx20800, nx20816, nx20830, nx20848, nx20862, nx20878, 
      nx20892, nx20920, nx20950, nx20988, nx21002, nx21004, nx21008, nx21016, 
      nx21034, nx21046, nx21062, nx21076, nx18631, nx18641, nx18651, nx18661, 
      nx18667, nx18681, nx18691, nx18701, nx18711, nx18721, nx18731, nx18741, 
      nx18751, nx18761, nx18771, nx18781, nx18791, nx18801, nx18811, nx18821, 
      nx18831, nx18841, nx18851, nx18861, nx18871, nx18881, nx18891, nx18901, 
      nx18911, nx18921, nx18931, nx18941, nx18951, nx18961, nx18971, nx18981, 
      nx18991, nx19001, nx19011, nx19021, nx19031, nx19041, nx19051, nx19061, 
      nx19071, nx19081, nx19091, nx19101, nx19111, nx19121, nx19131, nx19141, 
      nx19151, nx19161, nx19171, nx19181, nx19191, nx19201, nx19211, nx19221, 
      nx19231, nx19241, nx19251, nx19261, nx19271, nx19281, nx19291, nx19301, 
      nx19311, nx19321, nx19331, nx19341, nx19351, nx19361, nx19371, nx19381, 
      nx19391, nx19401, nx19411, nx19421, nx19431, nx19441, nx19451, nx19461, 
      nx19471, nx19481, nx19491, nx19501, nx19511, nx19521, nx19531, nx19541, 
      nx19551, nx19561, nx19571, nx19581, nx19591, nx19601, nx19611, nx19621, 
      nx19631, nx19641, nx19651, nx19661, nx19671, nx19681, nx19691, nx19701, 
      nx19711, nx19721, nx19731, nx19741, nx19751, nx19761, nx19771, nx19781, 
      nx19791, nx19801, nx19811, nx19821, nx19831, nx19841, nx19851, nx19861, 
      nx19871, nx19881, nx19891, nx19901, nx19911, nx19921, nx19931, nx19941, 
      nx19951, nx19961, nx19971, nx19981, nx19991, nx20001, nx20011, nx20021, 
      nx20031, nx20041, nx20051, nx20061, nx20071, nx20081, nx20091, nx20101, 
      nx20111, nx20121, nx20127, nx20141, nx20151, nx20161, nx20171, nx20181, 
      nx20191, nx20201, nx20211, nx20221, nx20231, nx20241, nx20251, nx20261, 
      nx20271, nx20281, nx20291, nx20301, nx20311, nx20321, nx20331, nx20341, 
      nx20351, nx20361, nx20371, nx20381, nx20391, nx20401, nx20411, nx20421, 
      nx20431, nx20441, nx20451, nx20461, nx20471, nx20481, nx20491, nx20501, 
      nx20511, nx20521, nx20531, nx20541, nx20551, nx20561, nx20571, nx20581, 
      nx20591, nx20601, nx20611, nx20621, nx20631, nx20641, nx20651, nx20661, 
      nx20671, nx20681, nx20691, nx20701, nx20711, nx20721, nx20731, nx20741, 
      nx20751, nx20761, nx20771, nx20781, nx20791, nx20801, nx20811, nx20821, 
      nx20831, nx20841, nx20851, nx20857, nx20871, nx20881, nx20891, nx20901, 
      nx20911, nx20921, nx20931, nx20941, nx20951, nx20961, nx20971, nx20981, 
      nx20991, nx21001, nx21011, nx21021, nx21031, nx21041, nx21051, nx21061, 
      nx21071, nx21081, nx21091, nx21101, nx21111, nx21121, nx21131, nx21141, 
      nx21151, nx21161, nx21171, nx21181, nx21191, nx21201, nx21211, nx21221, 
      nx21231, nx21241, nx21251, nx21261, nx21271, nx21281, nx21291, nx21301, 
      nx21311, nx21321, nx21331, nx21341, nx21351, nx21361, nx21371, nx21381, 
      nx21391, nx21401, nx21411, nx21421, nx21427, nx21441, nx21451, nx21461, 
      nx21471, nx21481, nx21491, nx21501, nx21511, nx21521, nx21531, nx21541, 
      nx21551, nx21561, nx21571, nx21581, nx21591, nx21601, nx21611, nx21621, 
      nx21631, nx21641, nx21651, nx21661, nx21671, nx21681, nx21691, nx21701, 
      nx21711, nx21721, nx21731, nx21741, nx21751, nx21761, nx21771, nx21781, 
      nx21791, nx21801, nx21811, nx21821, nx21831, nx21841, nx21851, nx21861, 
      nx21871, nx21881, nx21891, nx21901, nx21911, nx21921, nx21931, nx21941, 
      nx21951, nx21961, nx21971, nx21981, nx21991, nx22001, nx22011, nx22021, 
      nx22031, nx22041, nx22051, nx22061, nx22071, nx22081, nx22091, nx22101, 
      nx22111, nx22121, nx22131, nx22141, nx22151, nx22161, nx22171, nx22181, 
      nx22191, nx22201, nx22211, nx22221, nx22231, nx22241, nx22251, nx22261, 
      nx22271, nx22281, nx22291, nx22301, nx22311, nx22321, nx22331, nx22341, 
      nx22351, nx22361, nx22371, nx22381, nx22391, nx22401, nx22411, nx22421, 
      nx22431, nx22441, nx22451, nx22461, nx22471, nx22481, nx22491, nx22501, 
      nx22511, nx22521, nx22531, nx22541, nx22551, nx22561, nx22571, nx22581, 
      nx22591, nx22601, nx22611, nx22621, nx22631, nx22641, nx22651, nx22661, 
      nx22671, nx22681, nx22691, nx22701, nx22711, nx22721, nx22731, nx22741, 
      nx22751, nx22761, nx22771, nx22781, nx22791, nx22801, nx22811, nx22821, 
      nx22831, nx22841, nx22851, nx22861, nx22871, nx22881, nx22891, nx22901, 
      nx22907, nx22921, nx22931, nx22941, nx22951, nx22961, nx22971, nx22981, 
      nx22991, nx23001, nx23011, nx23021, nx23031, nx23041, nx23051, nx23061, 
      nx23071, nx23081, nx23091, nx23101, nx23111, nx23121, nx23131, nx23141, 
      nx23151, nx23161, nx23171, nx23181, nx23191, nx23201, nx23211, nx23221, 
      nx23231, nx23241, nx23251, nx23261, nx23271, nx23281, nx23291, nx23301, 
      nx23311, nx23321, nx23331, nx23341, nx23351, nx23361, nx23371, nx23381, 
      nx23391, nx23401, nx23411, nx23421, nx23431, nx23441, nx23451, nx23461, 
      nx23471, nx23481, nx23491, nx23501, nx23511, nx23521, nx23531, nx23541, 
      nx23551, nx23561, nx23571, nx23581, nx23591, nx23601, nx23611, nx23621, 
      nx23631, nx23641, nx23651, nx23661, nx23671, nx23681, nx23691, nx23701, 
      nx23711, nx23721, nx23731, nx23737, nx23751, nx23761, nx23771, nx23781, 
      nx23791, nx23801, nx23811, nx23821, nx23831, nx23841, nx23851, nx23861, 
      nx23871, nx23881, nx23891, nx23901, nx23911, nx23921, nx23931, nx23941, 
      nx23951, nx23961, nx23971, nx23981, nx23991, nx24001, nx24011, nx24021, 
      nx24031, nx24041, nx24051, nx24061, nx24071, nx24081, nx24091, nx24101, 
      nx24111, nx24121, nx24131, nx24141, nx24151, nx24161, nx24171, nx24181, 
      nx24191, nx24201, nx24211, nx24221, nx24231, nx24241, nx24251, nx24261, 
      nx24271, nx24281, nx24291, nx24301, nx24311, nx24321, nx24331, nx24341, 
      nx24351, nx24361, nx24371, nx24381, nx24391, nx24401, nx24411, nx24421, 
      nx24431, nx24441, nx24451, nx24461, nx24471, nx24481, nx24491, nx24501, 
      nx24511, nx24521, nx24531, nx24541, nx24551, nx24561, nx24567, nx24581, 
      nx24591, nx24601, nx24611, nx24621, nx24631, nx24641, nx24651, nx24661, 
      nx24671, nx24681, nx24691, nx24701, nx24711, nx24721, nx24731, nx24741, 
      nx24751, nx24761, nx24771, nx24781, nx24791, nx24801, nx24811, nx24821, 
      nx24831, nx24841, nx24851, nx24861, nx24871, nx24881, nx24891, nx24901, 
      nx24911, nx24921, nx24931, nx24941, nx24951, nx24961, nx24971, nx24981, 
      nx24991, nx25001, nx25011, nx25021, nx25031, nx25041, nx25051, nx25061, 
      nx25071, nx25081, nx25091, nx25101, nx25111, nx25121, nx25131, nx25141, 
      nx25151, nx25161, nx25171, nx25181, nx25191, nx25201, nx25211, nx25221, 
      nx25231, nx25241, nx25251, nx25261, nx25271, nx25281, nx25291, nx25301, 
      nx25311, nx25321, nx25331, nx25341, nx25351, nx25361, nx25371, nx25381, 
      nx25391, nx25401, nx25407, nx25421, nx25431, nx25441, nx25451, nx25461, 
      nx25471, nx25481, nx25491, nx25501, nx25511, nx25521, nx25531, nx25541, 
      nx25551, nx25561, nx25571, nx25581, nx25591, nx25601, nx25611, nx25621, 
      nx25631, nx25641, nx25651, nx25661, nx25671, nx25681, nx25691, nx25701, 
      nx25711, nx25721, nx25731, nx25741, nx25751, nx25761, nx25771, nx25781, 
      nx25791, nx25801, nx25811, nx25821, nx25831, nx25841, nx25851, nx25861, 
      nx25871, nx25881, nx25891, nx25901, nx25911, nx25921, nx25931, nx25941, 
      nx25951, nx25961, nx25971, nx25981, nx25991, nx26001, nx26011, nx26021, 
      nx26031, nx26041, nx26051, nx26061, nx26071, nx26081, nx26091, nx26101, 
      nx26111, nx26121, nx26131, nx26141, nx26151, nx26161, nx26171, nx26181, 
      nx26191, nx26201, nx26211, nx26221, nx26231, nx26241, nx26251, nx26261, 
      nx26271, nx26281, nx26291, nx26301, nx26311, nx26321, nx26331, nx26341, 
      nx26351, nx26361, nx26371, nx26381, nx26391, nx26401, nx26411, nx26421, 
      nx26431, nx26441, nx26451, nx26461, nx26471, nx26481, nx26491, nx26501, 
      nx26511, nx26521, nx26531, nx26541, nx26551, nx26561, nx26571, nx26581, 
      nx26591, nx26601, nx26607, nx26621, nx26631, nx26641, nx26651, nx26661, 
      nx26671, nx26681, nx26691, nx26701, nx26711, nx26721, nx26731, nx26741, 
      nx26751, nx26761, nx26771, nx26781, nx26791, nx26801, nx26811, nx26821, 
      nx26831, nx26841, nx26851, nx26861, nx26871, nx26881, nx26891, nx26901, 
      nx26911, nx26921, nx26931, nx26941, nx26951, nx26961, nx26971, nx26981, 
      nx26991, nx27001, nx27011, nx27021, nx27031, nx27041, nx27051, nx27061, 
      nx27071, nx27081, nx27091, nx27101, nx27111, nx27121, nx27131, nx27141, 
      nx27151, nx27161, nx27171, nx27181, nx27191, nx27201, nx27211, nx27221, 
      nx27231, nx27241, nx27251, nx27261, nx27271, nx27281, nx27291, nx27301, 
      nx27311, nx27321, nx27331, nx27341, nx27351, nx27361, nx27371, nx27381, 
      nx27391, nx27401, nx27411, nx27421, nx27431, nx27437, nx27451, nx27461, 
      nx27471, nx27481, nx27491, nx27501, nx27511, nx27521, nx27531, nx27541, 
      nx27551, nx27561, nx27571, nx27581, nx27591, nx27601, nx27611, nx27621, 
      nx27631, nx27641, nx27651, nx27661, nx27671, nx27681, nx27691, nx27701, 
      nx27711, nx27721, nx27731, nx27741, nx27751, nx27761, nx27771, nx27781, 
      nx27791, nx27801, nx27811, nx27821, nx27831, nx27841, nx27851, nx27861, 
      nx27871, nx27881, nx27891, nx27901, nx27911, nx27921, nx27931, nx27941, 
      nx27951, nx27961, nx27971, nx27981, nx27991, nx28001, nx28011, nx28021, 
      nx28031, nx28041, nx28051, nx28061, nx28071, nx28081, nx28091, nx28101, 
      nx28111, nx28121, nx28131, nx28141, nx28151, nx28161, nx28171, nx28181, 
      nx28191, nx28201, nx28211, nx28221, nx28231, nx28241, nx28251, nx28261, 
      nx28271, nx28277, nx28291, nx28301, nx28311, nx28321, nx28331, nx28341, 
      nx28351, nx28361, nx28371, nx28381, nx28391, nx28401, nx28411, nx28421, 
      nx28431, nx28441, nx28451, nx28461, nx28471, nx28481, nx28491, nx28501, 
      nx28511, nx28521, nx28531, nx28541, nx28551, nx28561, nx28571, nx28581, 
      nx28591, nx28601, nx28611, nx28621, nx28631, nx28641, nx28651, nx28661, 
      nx28671, nx28681, nx28691, nx28701, nx28711, nx28721, nx28731, nx28741, 
      nx28751, nx28761, nx28771, nx28781, nx28791, nx28801, nx28811, nx28821, 
      nx28831, nx28841, nx28851, nx28861, nx28871, nx28881, nx28891, nx28901, 
      nx28911, nx28921, nx28931, nx28941, nx28951, nx28961, nx28971, nx28981, 
      nx28991, nx29001, nx29011, nx29021, nx29031, nx29041, nx29051, nx29061, 
      nx29071, nx29081, nx29091, nx29101, nx29111, nx29121, nx29131, nx29141, 
      nx29151, nx29161, nx29171, nx29181, nx29191, nx29201, nx29211, nx29221, 
      nx29231, nx29241, nx29251, nx29261, nx29271, nx29281, nx29291, nx29301, 
      nx29311, nx29321, nx29331, nx29341, nx29351, nx29361, nx29371, nx29381, 
      nx29391, nx29401, nx29411, nx29421, nx29431, nx29441, nx29451, nx29461, 
      nx29471, nx29481, nx29491, nx29501, nx29511, nx29521, nx29531, nx29541, 
      nx29551, nx29561, nx29571, nx29581, nx29591, nx29601, nx29611, nx29621, 
      nx29631, nx29641, nx29651, nx29661, nx29671, nx29681, nx29691, nx29701, 
      nx29711, nx29721, nx29731, nx29741, nx29751, nx29761, nx29771, nx29781, 
      nx29791, nx29801, nx29811, nx29821, nx29831, nx29841, nx29851, nx29861, 
      nx29871, nx29881, nx29891, nx29901, nx29911, nx29921, nx29931, nx29941, 
      nx29951, nx29961, nx29971, nx29981, nx29991, nx30001, nx30011, nx30021, 
      nx30031, nx30041, nx30051, nx30061, nx30071, nx30081, nx30091, nx30101, 
      nx30111, nx30121, nx30131, nx30141, nx30151, nx30161, nx30171, nx30181, 
      nx30191, nx30201, nx30211, nx30221, nx30231, nx30241, nx30251, nx30261, 
      nx30271, nx30281, nx30291, nx30301, nx30311, nx30321, nx30331, nx30341, 
      nx30351, nx30361, nx30371, nx30381, nx30391, nx30401, nx30411, nx30421, 
      nx30431, nx30441, nx30451, nx30461, nx30471, nx30481, nx30491, nx30501, 
      nx30511, nx30521, nx30531, nx30541, nx30551, nx30561, nx30571, nx30581, 
      nx30591, nx30601, nx30611, nx30621, nx30631, nx30641, nx30651, nx30661, 
      nx30671, nx30681, nx30691, nx30701, nx30711, nx30721, nx30731, nx30741, 
      nx30751, nx30761, nx30771, nx30781, nx30791, nx30801, nx30811, nx30821, 
      nx30831, nx30841, nx30851, nx30861, nx30871, nx30881, nx30891, nx30901, 
      nx30911, nx30921, nx30931, nx30941, nx30951, nx30961, nx30971, nx30981, 
      nx30991, nx31001, nx31011, nx31021, nx31031, nx31041, nx31051, nx31061, 
      nx31071, nx31081, nx31091, nx31101, nx31111, nx31121, nx31131, nx31141, 
      nx31151, nx31161, nx31171, nx31181, nx31191, nx31201, nx31211, nx31221, 
      nx31231, nx31241, nx31251, nx31261, nx31271, nx31281, nx31291, nx31301, 
      nx31311, nx31321, nx31331, nx31341, nx31351, nx31361, nx31371, nx31381, 
      nx31391, nx31401, nx31411, nx31421, nx31431, nx31441, nx31451, nx31461, 
      nx31471, nx31481, nx31491, nx31501, nx31511, nx31521, nx31531, nx31541, 
      nx31551, nx31561, nx31571, nx31581, nx31591, nx31601, nx31611, nx31621, 
      nx31631, nx31641, nx31651, nx31661, nx31671, nx31681, nx31691, nx31701, 
      nx31711, nx31721, nx31731, nx31741, nx31751, nx31761, nx31771, nx31781, 
      nx31791, nx31801, nx31811, nx31821, nx31831, nx31841, nx31851, nx31861, 
      nx31871, nx31881, nx31896, nx31899, nx31906, nx31909, nx31914, nx31919, 
      nx31926, nx31930, nx31933, nx31938, nx31946, nx31948, nx31955, nx31957, 
      nx31959, nx31961, nx31966, nx31968, nx31970, nx31972, nx31974, nx31978, 
      nx31985, nx31991, nx32062, nx32072, nx32085, nx32089, nx32101, nx32103, 
      nx32113, nx32119, nx32126, nx32131, nx32137, nx32142, nx32144, nx32148, 
      nx32150, nx32164, nx32166, nx32175, nx32185, nx32197, nx32202, nx32208, 
      nx32212, nx32228, nx32230, nx32238, nx32246, nx32248, nx32251, nx32261, 
      nx32273, nx32274, nx32283, nx32287, nx32303, nx32305, nx32313, nx32321, 
      nx32323, nx32326, nx32336, nx32348, nx32349, nx32357, nx32361, nx32377, 
      nx32379, nx32387, nx32395, nx32397, nx32400, nx32410, nx32422, nx32423, 
      nx32432, nx32436, nx32452, nx32454, nx32462, nx32470, nx32472, nx32475, 
      nx32485, nx32497, nx32498, nx32506, nx32510, nx32526, nx32528, nx32536, 
      nx32544, nx32546, nx32549, nx32559, nx32571, nx32572, nx32581, nx32585, 
      nx32601, nx32603, nx32611, nx32619, nx32621, nx32624, nx32634, nx32646, 
      nx32647, nx32655, nx32659, nx32676, nx32678, nx32686, nx32689, nx32693, 
      nx32696, nx32700, nx32705, nx32709, nx32711, nx32714, nx32729, nx32733, 
      nx32744, nx32755, nx32766, nx32777, nx32788, nx32799, nx32810, nx32816, 
      nx32820, nx32833, nx32838, nx32886, nx32907, nx32912, nx32914, nx32999, 
      nx33001, nx33005, nx33011, nx33013, nx33016, nx33023, nx33026, nx33031, 
      nx33033, nx33037, nx33039, nx33042, nx33044, nx33048, nx33050, nx33053, 
      nx33056, nx33059, nx33067, nx33070, nx33072, nx33075, nx33077, nx33079, 
      nx33084, nx33086, nx33089, nx33101, nx33104, nx33106, nx33109, nx33111, 
      nx33113, nx33118, nx33120, nx33123, nx33135, nx33138, nx33140, nx33143, 
      nx33145, nx33147, nx33152, nx33154, nx33157, nx33169, nx33172, nx33174, 
      nx33177, nx33179, nx33181, nx33186, nx33188, nx33191, nx33203, nx33206, 
      nx33208, nx33211, nx33213, nx33215, nx33220, nx33222, nx33225, nx33236, 
      nx33238, nx33242, nx33244, nx33247, nx33249, nx33251, nx33254, nx33256, 
      nx33258, nx33261, nx33264, nx33267, nx33270, nx33273, nx33276, nx33280, 
      nx33289, nx33299, nx33302, nx33304, nx33312, nx33315, nx33325, nx33326, 
      nx33330, nx33340, nx33341, nx33345, nx33355, nx33356, nx33360, nx33370, 
      nx33371, nx33375, nx33385, nx33386, nx33390, nx33400, nx33401, nx33405, 
      nx33415, nx33416, nx33421, nx33429, nx33432, nx33436, nx33444, nx33447, 
      nx33450, nx33453, nx33463, nx33474, nx33485, nx33496, nx33507, nx33518, 
      nx33529, nx33540, nx33546, nx33550, nx33563, nx33610, nx33631, nx33636, 
      nx33638, nx33687, nx33689, nx33693, nx33699, nx33701, nx33704, nx33709, 
      nx33714, nx33719, nx33721, nx33725, nx33727, nx33730, nx33734, nx33738, 
      nx33740, nx33743, nx33746, nx33749, nx33757, nx33760, nx33762, nx33765, 
      nx33767, nx33769, nx33771, nx33776, nx33778, nx33781, nx33793, nx33796, 
      nx33798, nx33801, nx33803, nx33805, nx33807, nx33812, nx33814, nx33817, 
      nx33829, nx33832, nx33834, nx33837, nx33839, nx33841, nx33843, nx33848, 
      nx33850, nx33853, nx33865, nx33868, nx33870, nx33873, nx33875, nx33877, 
      nx33879, nx33884, nx33886, nx33889, nx33901, nx33904, nx33906, nx33909, 
      nx33911, nx33913, nx33915, nx33920, nx33922, nx33925, nx33936, nx33938, 
      nx33942, nx33944, nx33947, nx33949, nx33951, nx33953, nx33956, nx33958, 
      nx33960, nx33963, nx33966, nx33969, nx33972, nx33975, nx33978, nx33982, 
      nx33985, nx33989, nx33999, nx34000, nx34004, nx34014, nx34015, nx34019, 
      nx34029, nx34030, nx34034, nx34044, nx34045, nx34049, nx34059, nx34060, 
      nx34064, nx34074, nx34075, nx34079, nx34089, nx34090, nx34095, nx34097, 
      nx34114, nx34125, nx34128, nx34139, nx34150, nx34161, nx34172, nx34183, 
      nx34194, nx34205, nx34211, nx34215, nx34228, nx34275, nx34296, nx34301, 
      nx34303, nx34352, nx34354, nx34358, nx34364, nx34366, nx34369, nx34374, 
      nx34379, nx34384, nx34386, nx34390, nx34392, nx34395, nx34399, nx34403, 
      nx34405, nx34408, nx34411, nx34414, nx34422, nx34425, nx34427, nx34430, 
      nx34432, nx34434, nx34436, nx34441, nx34443, nx34446, nx34458, nx34461, 
      nx34463, nx34466, nx34468, nx34470, nx34472, nx34477, nx34479, nx34482, 
      nx34494, nx34497, nx34499, nx34502, nx34504, nx34506, nx34508, nx34513, 
      nx34515, nx34518, nx34530, nx34533, nx34535, nx34538, nx34540, nx34542, 
      nx34544, nx34549, nx34551, nx34554, nx34566, nx34569, nx34571, nx34574, 
      nx34576, nx34578, nx34580, nx34585, nx34587, nx34590, nx34601, nx34603, 
      nx34607, nx34609, nx34612, nx34614, nx34616, nx34618, nx34621, nx34623, 
      nx34625, nx34628, nx34631, nx34634, nx34637, nx34640, nx34643, nx34647, 
      nx34650, nx34654, nx34664, nx34665, nx34669, nx34679, nx34680, nx34684, 
      nx34694, nx34695, nx34699, nx34709, nx34710, nx34714, nx34724, nx34725, 
      nx34729, nx34739, nx34740, nx34744, nx34754, nx34755, nx34760, nx34762, 
      nx34765, nx34769, nx34773, nx34775, nx34777, nx34780, nx34782, nx34784, 
      nx34787, nx34791, nx34793, nx34797, nx34801, nx34803, nx34805, nx34808, 
      nx34810, nx34812, nx34815, nx34819, nx34821, nx34825, nx34829, nx34831, 
      nx34833, nx34836, nx34838, nx34840, nx34843, nx34847, nx34849, nx34853, 
      nx34857, nx34859, nx34861, nx34864, nx34866, nx34868, nx34871, nx34875, 
      nx34877, nx34881, nx34885, nx34887, nx34889, nx34892, nx34894, nx34896, 
      nx34899, nx34903, nx34905, nx34909, nx34913, nx34915, nx34917, nx34920, 
      nx34922, nx34924, nx34927, nx34931, nx34933, nx34939, nx34941, nx34943, 
      nx34946, nx34948, nx34950, nx34953, nx34957, nx34959, nx34965, nx34967, 
      nx34971, nx34973, nx34983, nx34987, nx34993, nx35009, nx35020, nx35031, 
      nx35042, nx35053, nx35064, nx35075, nx35081, nx35085, nx35098, nx35145, 
      nx35166, nx35171, nx35173, nx35222, nx35224, nx35228, nx35234, nx35236, 
      nx35239, nx35244, nx35249, nx35254, nx35256, nx35260, nx35262, nx35265, 
      nx35269, nx35273, nx35275, nx35278, nx35281, nx35284, nx35292, nx35295, 
      nx35297, nx35300, nx35302, nx35304, nx35306, nx35311, nx35313, nx35316, 
      nx35328, nx35331, nx35333, nx35336, nx35338, nx35340, nx35342, nx35347, 
      nx35349, nx35352, nx35364, nx35367, nx35369, nx35372, nx35374, nx35376, 
      nx35378, nx35383, nx35385, nx35388, nx35400, nx35403, nx35405, nx35408, 
      nx35410, nx35412, nx35414, nx35419, nx35421, nx35424, nx35436, nx35439, 
      nx35441, nx35444, nx35446, nx35448, nx35450, nx35455, nx35457, nx35460, 
      nx35471, nx35473, nx35477, nx35479, nx35482, nx35484, nx35486, nx35488, 
      nx35491, nx35493, nx35495, nx35498, nx35501, nx35504, nx35507, nx35510, 
      nx35513, nx35517, nx35520, nx35524, nx35534, nx35535, nx35539, nx35549, 
      nx35550, nx35554, nx35564, nx35565, nx35569, nx35579, nx35580, nx35584, 
      nx35594, nx35595, nx35599, nx35609, nx35610, nx35614, nx35624, nx35625, 
      nx35633, nx35635, nx35647, nx35658, nx35669, nx35680, nx35691, nx35702, 
      nx35713, nx35719, nx35723, nx35736, nx35783, nx35804, nx35809, nx35811, 
      nx35860, nx35862, nx35866, nx35872, nx35874, nx35877, nx35882, nx35887, 
      nx35892, nx35894, nx35898, nx35900, nx35903, nx35907, nx35911, nx35913, 
      nx35916, nx35919, nx35922, nx35930, nx35933, nx35935, nx35938, nx35940, 
      nx35942, nx35944, nx35949, nx35951, nx35954, nx35966, nx35969, nx35971, 
      nx35974, nx35976, nx35978, nx35980, nx35985, nx35987, nx35990, nx36002, 
      nx36005, nx36007, nx36010, nx36012, nx36014, nx36016, nx36021, nx36023, 
      nx36026, nx36038, nx36041, nx36043, nx36046, nx36048, nx36050, nx36052, 
      nx36057, nx36059, nx36062, nx36074, nx36077, nx36079, nx36082, nx36084, 
      nx36086, nx36088, nx36093, nx36095, nx36098, nx36109, nx36111, nx36115, 
      nx36117, nx36120, nx36122, nx36124, nx36126, nx36129, nx36131, nx36133, 
      nx36136, nx36139, nx36142, nx36145, nx36148, nx36151, nx36155, nx36158, 
      nx36162, nx36172, nx36173, nx36177, nx36187, nx36188, nx36192, nx36202, 
      nx36203, nx36207, nx36217, nx36218, nx36222, nx36232, nx36233, nx36237, 
      nx36247, nx36248, nx36252, nx36262, nx36263, nx36271, nx36273, nx36284, 
      nx36295, nx36306, nx36317, nx36328, nx36339, nx36350, nx36356, nx36360, 
      nx36373, nx36420, nx36441, nx36446, nx36448, nx36497, nx36499, nx36503, 
      nx36509, nx36511, nx36514, nx36519, nx36524, nx36529, nx36531, nx36535, 
      nx36537, nx36540, nx36544, nx36548, nx36550, nx36553, nx36556, nx36559, 
      nx36567, nx36570, nx36572, nx36575, nx36577, nx36579, nx36581, nx36586, 
      nx36588, nx36591, nx36603, nx36606, nx36608, nx36611, nx36613, nx36615, 
      nx36617, nx36622, nx36624, nx36627, nx36639, nx36642, nx36644, nx36647, 
      nx36649, nx36651, nx36653, nx36658, nx36660, nx36663, nx36675, nx36678, 
      nx36680, nx36683, nx36685, nx36687, nx36689, nx36694, nx36696, nx36699, 
      nx36711, nx36714, nx36716, nx36719, nx36721, nx36723, nx36725, nx36730, 
      nx36732, nx36735, nx36746, nx36748, nx36752, nx36754, nx36757, nx36759, 
      nx36761, nx36763, nx36766, nx36768, nx36770, nx36773, nx36776, nx36779, 
      nx36782, nx36785, nx36788, nx36792, nx36795, nx36799, nx36809, nx36810, 
      nx36814, nx36824, nx36825, nx36829, nx36839, nx36840, nx36844, nx36854, 
      nx36855, nx36859, nx36869, nx36870, nx36874, nx36884, nx36885, nx36889, 
      nx36899, nx36900, nx36903, nx36907, nx36909, nx36920, nx36931, nx36942, 
      nx36953, nx36964, nx36975, nx36986, nx36992, nx36996, nx37009, nx37056, 
      nx37077, nx37082, nx37084, nx37133, nx37135, nx37139, nx37145, nx37147, 
      nx37150, nx37155, nx37160, nx37165, nx37167, nx37171, nx37173, nx37176, 
      nx37180, nx37184, nx37186, nx37189, nx37192, nx37195, nx37203, nx37206, 
      nx37208, nx37211, nx37213, nx37215, nx37217, nx37222, nx37224, nx37227, 
      nx37239, nx37242, nx37244, nx37247, nx37249, nx37251, nx37253, nx37258, 
      nx37260, nx37263, nx37275, nx37278, nx37280, nx37283, nx37285, nx37287, 
      nx37289, nx37294, nx37296, nx37299, nx37311, nx37314, nx37316, nx37319, 
      nx37321, nx37323, nx37325, nx37330, nx37332, nx37335, nx37347, nx37350, 
      nx37352, nx37355, nx37357, nx37359, nx37361, nx37366, nx37368, nx37371, 
      nx37382, nx37384, nx37388, nx37390, nx37393, nx37395, nx37397, nx37399, 
      nx37402, nx37404, nx37406, nx37409, nx37412, nx37415, nx37418, nx37421, 
      nx37424, nx37428, nx37431, nx37435, nx37445, nx37446, nx37450, nx37460, 
      nx37461, nx37465, nx37475, nx37476, nx37480, nx37490, nx37491, nx37495, 
      nx37505, nx37506, nx37510, nx37520, nx37521, nx37525, nx37535, nx37536, 
      nx37540, nx37544, nx37548, nx37550, nx37552, nx37555, nx37557, nx37559, 
      nx37562, nx37566, nx37568, nx37572, nx37576, nx37578, nx37580, nx37583, 
      nx37585, nx37587, nx37590, nx37594, nx37596, nx37600, nx37604, nx37606, 
      nx37608, nx37611, nx37613, nx37615, nx37618, nx37622, nx37624, nx37628, 
      nx37632, nx37634, nx37636, nx37639, nx37641, nx37643, nx37646, nx37650, 
      nx37652, nx37656, nx37660, nx37662, nx37664, nx37667, nx37669, nx37671, 
      nx37674, nx37678, nx37680, nx37684, nx37688, nx37690, nx37692, nx37695, 
      nx37697, nx37699, nx37702, nx37706, nx37708, nx37714, nx37716, nx37718, 
      nx37721, nx37723, nx37725, nx37728, nx37732, nx37734, nx37740, nx37742, 
      nx37752, nx37756, nx37760, nx37762, nx37772, nx37776, nx37785, nx37787, 
      nx37799, nx37810, nx37821, nx37832, nx37843, nx37854, nx37865, nx37871, 
      nx37875, nx37888, nx37935, nx37956, nx37961, nx37963, nx38012, nx38014, 
      nx38018, nx38024, nx38026, nx38029, nx38034, nx38039, nx38044, nx38046, 
      nx38050, nx38052, nx38055, nx38059, nx38063, nx38065, nx38068, nx38071, 
      nx38074, nx38082, nx38085, nx38087, nx38090, nx38092, nx38094, nx38096, 
      nx38101, nx38103, nx38106, nx38118, nx38121, nx38123, nx38126, nx38128, 
      nx38130, nx38132, nx38137, nx38139, nx38142, nx38154, nx38157, nx38159, 
      nx38162, nx38164, nx38166, nx38168, nx38173, nx38175, nx38178, nx38190, 
      nx38193, nx38195, nx38198, nx38200, nx38202, nx38204, nx38209, nx38211, 
      nx38214, nx38226, nx38229, nx38231, nx38234, nx38236, nx38238, nx38240, 
      nx38245, nx38247, nx38250, nx38261, nx38263, nx38267, nx38269, nx38272, 
      nx38274, nx38276, nx38278, nx38281, nx38283, nx38285, nx38288, nx38291, 
      nx38294, nx38297, nx38300, nx38303, nx38307, nx38310, nx38314, nx38324, 
      nx38325, nx38329, nx38339, nx38340, nx38344, nx38354, nx38355, nx38359, 
      nx38369, nx38370, nx38374, nx38384, nx38385, nx38389, nx38399, nx38400, 
      nx38404, nx38414, nx38415, nx38423, nx38425, nx38436, nx38447, nx38458, 
      nx38469, nx38480, nx38491, nx38502, nx38508, nx38512, nx38525, nx38572, 
      nx38593, nx38598, nx38600, nx38649, nx38651, nx38655, nx38661, nx38663, 
      nx38666, nx38671, nx38676, nx38681, nx38683, nx38687, nx38689, nx38692, 
      nx38696, nx38700, nx38702, nx38705, nx38708, nx38711, nx38719, nx38722, 
      nx38724, nx38727, nx38729, nx38731, nx38733, nx38738, nx38740, nx38743, 
      nx38755, nx38758, nx38760, nx38763, nx38765, nx38767, nx38769, nx38774, 
      nx38776, nx38779, nx38791, nx38794, nx38796, nx38799, nx38801, nx38803, 
      nx38805, nx38810, nx38812, nx38815, nx38827, nx38830, nx38832, nx38835, 
      nx38837, nx38839, nx38841, nx38846, nx38848, nx38851, nx38863, nx38866, 
      nx38868, nx38871, nx38873, nx38875, nx38877, nx38882, nx38884, nx38887, 
      nx38898, nx38900, nx38904, nx38906, nx38909, nx38911, nx38913, nx38915, 
      nx38918, nx38920, nx38922, nx38925, nx38928, nx38931, nx38934, nx38937, 
      nx38940, nx38944, nx38947, nx38951, nx38961, nx38962, nx38966, nx38976, 
      nx38977, nx38981, nx38991, nx38992, nx38996, nx39006, nx39007, nx39011, 
      nx39021, nx39022, nx39026, nx39036, nx39037, nx39041, nx39051, nx39052, 
      nx39057, nx39059, nx39070, nx39081, nx39092, nx39103, nx39114, nx39125, 
      nx39136, nx39142, nx39146, nx39159, nx39206, nx39227, nx39232, nx39234, 
      nx39283, nx39285, nx39289, nx39295, nx39297, nx39300, nx39305, nx39310, 
      nx39315, nx39317, nx39321, nx39323, nx39326, nx39330, nx39334, nx39336, 
      nx39339, nx39342, nx39345, nx39353, nx39356, nx39358, nx39361, nx39363, 
      nx39365, nx39367, nx39372, nx39374, nx39377, nx39389, nx39392, nx39394, 
      nx39397, nx39399, nx39401, nx39403, nx39408, nx39410, nx39413, nx39425, 
      nx39428, nx39430, nx39433, nx39435, nx39437, nx39439, nx39444, nx39446, 
      nx39449, nx39461, nx39464, nx39466, nx39469, nx39471, nx39473, nx39475, 
      nx39480, nx39482, nx39485, nx39497, nx39500, nx39502, nx39505, nx39507, 
      nx39509, nx39511, nx39516, nx39518, nx39521, nx39532, nx39534, nx39538, 
      nx39540, nx39543, nx39545, nx39547, nx39549, nx39552, nx39554, nx39556, 
      nx39559, nx39562, nx39565, nx39568, nx39571, nx39574, nx39578, nx39581, 
      nx39585, nx39595, nx39596, nx39600, nx39610, nx39611, nx39615, nx39625, 
      nx39626, nx39630, nx39640, nx39641, nx39645, nx39655, nx39656, nx39660, 
      nx39670, nx39671, nx39675, nx39685, nx39686, nx39690, nx39694, nx39698, 
      nx39700, nx39702, nx39705, nx39707, nx39709, nx39712, nx39716, nx39718, 
      nx39722, nx39726, nx39728, nx39730, nx39733, nx39735, nx39737, nx39740, 
      nx39744, nx39746, nx39750, nx39754, nx39756, nx39758, nx39761, nx39763, 
      nx39765, nx39768, nx39772, nx39774, nx39778, nx39782, nx39784, nx39786, 
      nx39789, nx39791, nx39793, nx39796, nx39800, nx39802, nx39806, nx39810, 
      nx39812, nx39814, nx39817, nx39819, nx39821, nx39824, nx39828, nx39830, 
      nx39834, nx39838, nx39840, nx39842, nx39845, nx39847, nx39849, nx39852, 
      nx39856, nx39858, nx39864, nx39866, nx39868, nx39871, nx39873, nx39875, 
      nx39878, nx39882, nx39884, nx39890, nx39892, nx39902, nx39906, nx39910, 
      nx39912, nx39922, nx39926, nx39930, nx39934, nx39938, nx39940, nx39947, 
      nx39950, nx39957, nx39959, nx39962, nx39971, nx39973, nx39982, nx39986, 
      nx39988, nx39995, nx39998, nx40005, nx40007, nx40010, nx40019, nx40021, 
      nx40030, nx40034, nx40036, nx40043, nx40046, nx40053, nx40055, nx40058, 
      nx40067, nx40069, nx40078, nx40082, nx40084, nx40091, nx40094, nx40101, 
      nx40103, nx40106, nx40115, nx40117, nx40126, nx40130, nx40132, nx40139, 
      nx40142, nx40149, nx40151, nx40154, nx40163, nx40165, nx40174, nx40178, 
      nx40180, nx40187, nx40190, nx40197, nx40199, nx40202, nx40211, nx40213, 
      nx40224, nx40226, nx40233, nx40236, nx40243, nx40245, nx40248, nx40257, 
      nx40259, nx40270, nx40272, nx40283, nx40287, nx40295, nx40297, nx40308, 
      nx40312, nx40326, nx40328, nx40332, nx40364, nx40367, nx40369, nx40405, 
      nx40437, nx40440, nx40442, nx40478, nx40510, nx40513, nx40515, nx40551, 
      nx40583, nx40586, nx40588, nx40624, nx40656, nx40659, nx40661, nx40697, 
      nx40729, nx40732, nx40734, nx40800, nx40803, nx40805, nx40853, nx40857, 
      nx40874, nx40879, nx40885, nx40890, nx40895, nx40900, nx40906, nx40911, 
      nx40916, nx40921, nx40927, nx40932, nx40937, nx40942, nx40947, nx40950, 
      nx40952, nx40954, nx40956, nx40959, nx40961, nx40963, nx40965, nx40968, 
      nx40970, nx40972, nx40974, nx40977, nx40979, nx40981, nx40983, nx40985, 
      nx40998, nx41000, nx41002, nx41005, nx41007, nx41009, nx41011, nx41014, 
      nx41016, nx41018, nx41020, nx41023, nx41025, nx41027, nx41029, nx41031, 
      nx41034, nx41036, nx41038, nx41040, nx41042, nx41044, nx41046, nx41048, 
      nx41050, nx41052, nx41054, nx41056, nx41058, nx41060, nx41062, nx41064, 
      nx41066, nx41068, nx41070, nx41072, nx41075, nx41077, nx41080, nx41082, 
      nx41084, nx41086, nx41089, nx41091, nx41093, nx41095, nx41098, nx41100, 
      nx41102, nx41104, nx41107, nx41109, nx41111, nx41113, nx41115, nx41118, 
      nx41120, nx41122, nx41124, nx41126, nx41128, nx41130, nx41132, nx41134, 
      nx41136, nx41138, nx41140, nx41142, nx41144, nx41146, nx41148, nx41150, 
      nx41152, nx41154, nx41156, nx41158, nx41161, nx41163, nx41165, nx41167, 
      nx41170, nx41172, nx41174, nx41176, nx41179, nx41181, nx41183, nx41185, 
      nx41188, nx41190, nx41192, nx41194, nx41198, nx41200, nx41202, nx41204, 
      nx41207, nx41209, nx41211, nx41213, nx41216, nx41218, nx41220, nx41222, 
      nx41225, nx41227, nx41229, nx41231, nx41233, nx41236, nx41238, nx41240, 
      nx41242, nx41245, nx41247, nx41249, nx41251, nx41254, nx41256, nx41258, 
      nx41260, nx41263, nx41265, nx41267, nx41269, nx41273, nx41275, nx41277, 
      nx41279, nx41282, nx41284, nx41286, nx41288, nx41291, nx41293, nx41295, 
      nx41297, nx41300, nx41302, nx41304, nx41306, nx41310, nx41313, nx41319, 
      nx41321, nx41325, nx41328, nx41330, nx41332, nx41348, nx41354, nx41357, 
      nx41360, nx41362, nx41371, nx41373, nx41375, nx41377, nx41379, nx41381, 
      nx41383, nx41385, nx41387, nx41389, nx41391, nx41397, nx41405, nx41407, 
      nx41409, nx41411, nx41413, nx41415, nx41417, nx41419, nx41421, nx41425, 
      nx41429, nx41435, nx41439, nx41443, nx41447, nx41453, nx41457, nx41461, 
      nx41469, nx41471, nx41473, nx41475, nx41477, nx41479, nx41481, nx41483, 
      nx41485, nx41487, nx41489, nx41491, nx41493, nx41495, nx41497, nx41499, 
      nx41501, nx41503, nx41505, nx41515, nx41521, nx41523, nx41525, nx41527, 
      nx41529, nx41531, nx41533, nx41535, nx41563, nx41565, nx41575, nx41577, 
      nx41579, nx41581, nx41583, nx41585, nx41587, nx41589, nx41591, nx41593, 
      nx41595, nx41597, nx41599, nx41601, nx41603, nx41605, nx41607, nx41609, 
      nx41611, nx41613, nx41615, nx41617, nx41619, nx41621, nx41623, nx41625, 
      nx41627, nx41629, nx41631, nx41633, nx41635, nx41637, nx41639, nx41641, 
      nx41643, nx41645, nx41647, nx41649, nx41651, nx41653, nx41655, nx41657, 
      nx41659, nx41661, nx41663, nx41665, nx41667, nx41669, nx41671, nx41673, 
      nx41675, nx41677, nx41679, nx41681, nx41683, nx41685, nx41687, nx41689, 
      nx41691, nx41693, nx41695, nx41697, nx41699, nx41701, nx41703, nx41705, 
      nx41707, nx41721, nx41729, nx41731, nx41733, nx41741, nx41743, nx41745, 
      nx41747, nx41749, nx41751, nx41753, nx41755, nx41757, nx41759, nx41761, 
      nx41763, nx41765, nx41767, nx41769, nx41771, nx41773, nx41775, nx41777, 
      nx41779, nx41781, nx41783, nx41785, nx41787, nx41789, nx41791, nx41793, 
      nx41795, nx41797, nx41799, nx41801, nx41803, nx41805, nx41807, nx41809, 
      nx41811, nx41813, nx41815, nx41817, nx41819, nx41821, nx41833, nx41847, 
      nx41855, nx41857, nx41859, nx41861, nx41863, nx41865, nx41879, nx41887, 
      nx41889, nx41891, nx41893, nx41895, nx41905, nx41919, nx41927, nx41929, 
      nx41931, nx41933, nx41935, nx41937, nx41951, nx41959, nx41961, nx41963, 
      nx41965, nx41967, nx41969, nx41983, nx41991, nx41993, nx41995, nx41997, 
      nx41999, nx42001, nx42015, nx42023, nx42025, nx42027, nx42029, nx42031, 
      nx42041, nx42055, nx42063, nx42065, nx42067, nx42069, nx42071, nx42073, 
      nx42087, nx42095, nx42097, nx42099, nx42101, nx42103, nx42105, nx42119, 
      nx42127, nx42129, nx42131, nx42133, nx42135, nx42161, nx42163, nx42165, 
      nx42167, nx42169, nx42171, nx42173, nx42175, nx42177, nx42179, nx42181, 
      nx42183, nx42185, nx42187, nx42189, nx42191, nx42193, nx42195, nx42197, 
      nx42199, nx42201, nx42203, nx42205, nx42207, nx42209, nx42211, nx42213, 
      nx42215, nx42217, nx42219, nx42227, nx42229, nx42231, nx42233, nx42235, 
      nx42237, nx42239, nx42241, nx42243, nx42245, nx42247, nx42249, nx42251, 
      nx42253, nx42255, nx42257, nx42259, nx42261, nx42263, nx42271, nx42273, 
      nx42277, nx42279, nx42281, nx42283, nx42285, nx42287, nx42289, nx42291, 
      nx42293, nx42295, nx42299, nx42301, nx42303, nx42311, nx42313, nx42315, 
      nx42317, nx42373, nx42375, nx42377, nx42379, nx42381, nx42383, nx42385, 
      nx42387, nx42389, nx42391, nx42393, nx42395, nx42397, nx42443, nx42445, 
      nx42447, nx42449, nx42451, nx42453, nx42455, nx42457, nx42459, nx42461, 
      nx42463, nx42465, nx42467, nx42469, nx42471, nx42473, nx42475, nx42477, 
      nx42479, nx42481, nx42483, nx42485, nx42497, nx42499, nx42501, nx42503, 
      nx42505, nx42507, nx42509, nx42511, nx42513, nx42515, nx42517, nx42519, 
      nx42521, nx42527, nx42529, nx42539, nx42541, nx42543, nx42545, nx42547, 
      nx42549, nx42551, nx42553, nx42555, nx42557, nx42559, nx42561, nx42563, 
      nx42565, nx42567, nx42569, nx42571, nx42573, nx42575, nx42577, nx42579, 
      nx42581, nx42583, nx42585, nx42587, nx42589, nx42591, nx42593, nx42595, 
      nx42597, nx42599, nx42601, nx42603, nx42605, nx42607, nx42609, nx42611, 
      nx42613, nx42615, nx42617, nx42619, nx42621, nx42623, nx42625, nx42627, 
      nx42631, nx42633, nx42635, nx42637, nx42639, nx42641, nx42643, nx42645, 
      nx42647, nx42651, nx42653, nx42655, nx42657, nx42659, nx42661, nx42663, 
      nx42665, nx42667, nx42669, nx42671, nx42673, nx42675, nx42677, nx42679, 
      nx42681, nx42683, nx42685, nx42687, nx42689, nx42697, nx42699, nx42701, 
      nx42703, nx42705, nx42707, nx42709, nx42711, nx42713, nx42715, nx42717, 
      nx42719, nx42721, nx42723, nx42725, nx42727, nx42729, nx42731, nx42733, 
      nx42735, nx42737, nx42739, nx42741, nx42743, nx42745, nx42747, nx42749, 
      nx42751, nx42753, nx42755, nx42757, nx42759, nx42761, nx42763, nx42765, 
      nx42767, nx42769, nx42771, nx42773, nx42775, nx42789, nx42791, nx42793, 
      nx42795, nx42797, nx42799, nx42801, nx42803, nx42805, nx42809, nx42811, 
      nx42813, nx42815, nx42817, nx42819, nx42825, nx42827, nx42829, nx42831, 
      nx42833, nx42835, nx42837, nx42839, nx42841, nx42843, nx42845, nx42847, 
      nx42849, nx42851, nx42853, nx42855, nx42857, nx42859, nx42861, nx42863, 
      nx42865, nx42867, nx42869, nx42871, nx42873, nx42875, nx42877, nx42879, 
      nx42881, nx42883, nx42885, nx42887, nx42889, nx42891, nx42893, nx42895, 
      nx42897, nx42899, nx42901, nx42903, nx42905, nx42907, nx42909, nx42911, 
      nx42913, nx42915, nx42917, nx42919, nx42921, nx42923, nx42925, nx42927, 
      nx42929, nx42931, nx42933, nx42935, nx42937, nx42939, nx42941, nx42943, 
      nx42945, nx42947, nx42949, nx42951, nx42953, nx42955, nx42957, nx42959, 
      nx42961, nx42963, nx42965, nx42967, nx42969, nx42971, nx42973, nx42975, 
      nx42977, nx42979, nx42981, nx42983, nx42985, nx42987, nx42989, nx42991, 
      nx42993, nx42995, nx42997, nx42999, nx43001, nx43003, nx43005, nx43007, 
      nx43009, nx43011, nx43013, nx43015, nx43017, nx43019, nx43021, nx43023, 
      nx43025, nx43027, nx43029, nx43031, nx43033, nx43035, nx43037, nx43039, 
      nx43041, nx43043, nx43045, nx43047, nx43049, nx43051, nx43053, nx43055, 
      nx43057, nx43059, nx43061, nx43063, nx43065, nx43067, nx43069, nx43071, 
      nx43073, nx43075, nx43077, nx43079, nx43081, nx43083, nx43085, nx43087, 
      nx43089, nx43091, nx43093, nx43095, nx43097, nx43099, nx43101, nx43103, 
      nx43105, nx43107, nx43109, nx43111, nx43113, nx43115, nx43117, nx43119, 
      nx43121, nx43123, nx43125, nx43127, nx43129, nx43131, nx43133, nx43135, 
      nx43137, nx43139, nx43141, nx43143, nx43145, nx43147, nx43149, nx43151, 
      nx43153, nx43155, nx43157, nx43159, nx43161, nx43163, nx43165, nx43167, 
      nx43169, nx43171, nx43173, nx43175, nx43177, nx43179, nx43181, nx43183, 
      nx43185, nx43187, nx43189, nx43191, nx43193, nx43195, nx43197, nx43199, 
      nx43201, nx43203, nx43205, nx43207, nx43209, nx43211, nx43213, nx43215, 
      nx43217, nx43219, nx43221, nx43223, nx43225, nx43227, nx43229, nx43231, 
      nx43233, nx43235, nx43237, nx43239, nx43241, nx43243, nx43245, nx43247, 
      nx43249, nx43251, nx43253, nx43255, nx43257, nx43259, nx43261, nx43263, 
      nx43265, nx43267, nx43269, nx43271, nx43273, nx43275, nx43277, nx43279, 
      nx43281, nx43283, nx43285, nx43287, nx43289, nx43291, nx43293, nx43295, 
      nx43297, nx43299, nx43301, nx43303, nx43305, nx43307, nx43309, nx43311, 
      nx43313, nx43315, nx43317, nx43319, nx43321, nx43323, nx43325, nx43327, 
      nx43329, nx43331, nx43333, nx43335, nx43337, nx43339, nx43341, nx43343, 
      nx43345, nx43347, nx43349, nx43351, nx43353, nx43355, nx43357, nx43359, 
      nx43361, nx43363, nx43365, nx43367, nx43369, nx43371, nx43373, nx43375, 
      nx43377, nx43379, nx43381, nx43383, nx43385, nx43387, nx43389, nx43391, 
      nx43393, nx43395, nx43397, nx43399, nx43401, nx43403, nx43405, nx43407, 
      nx43409, nx43411, nx43413, nx43415, nx43417, nx43419, nx43421, nx43423, 
      nx43425, nx43427, nx43429, nx43431, nx43433, nx43435, nx43437, nx43439, 
      nx43445, nx43447, nx43449, nx43451, nx43453, nx43455, nx43457, nx43459, 
      nx43461, nx43463, nx43465, nx43467, nx43469, nx43471, nx43473, nx43475, 
      nx43477, nx43479, nx43481, nx43483, nx43485, nx43487, nx43489, nx43491, 
      nx43493, nx43495, nx43497, nx43499, nx43501, nx43503, nx43505, nx43507, 
      nx43509, nx43511, nx43513, nx43515, nx43517, nx43519, nx43521: 
   std_logic ;

begin
   enable_read <= enable_read_EXMPLR ;
   answer(3) <= answer_3_EXMPLR ;
   answer(2) <= answer_2_EXMPLR ;
   answer(1) <= answer_1_EXMPLR ;
   answer(0) <= answer_0_EXMPLR ;
   ix17959 : fake_gnd port map ( Y=>initiate);
   max_calc_reg_done_comp : dffr port map ( Q=>done_comp, QB=>OPEN, D=>
      nx31831, CLK=>clk, R=>rst);
   ix31832 : or02 port map ( Y=>nx31831, A0=>done_comp, A1=>nx20950);
   ix20951 : nor04_2x port map ( Y=>nx20950, A0=>nx18189, A1=>nx31896, A2=>
      nx1782, A3=>nx18191);
   ix20082 : oai22 port map ( Y=>nx20081, A0=>nx31896, A1=>nx32700, B0=>
      nx43031, B1=>nx1714);
   max_calc_reg_start : dffr port map ( Q=>max_calc_start, QB=>nx31896, D=>
      nx20071, CLK=>clk, R=>rst);
   ix20072 : nand02 port map ( Y=>nx20071, A0=>nx31896, A1=>nx31899);
   ix31900 : nand02 port map ( Y=>nx31899, A0=>start_comp, A1=>nx31896);
   reg_start_comp : dffr port map ( Q=>start_comp, QB=>OPEN, D=>nx20061, CLK
      =>clk, R=>rst);
   ix20062 : or02 port map ( Y=>nx20061, A0=>start_comp, A1=>nx41381);
   ix20052 : oai22 port map ( Y=>nx20051, A0=>nx31909, A1=>nx32689, B0=>
      nx31906, B1=>nx42877);
   ix31910 : aoi221 port map ( Y=>nx31909, A0=>nx42259, A1=>nx18159, B0=>
      nx31961, B1=>nx41389, C0=>nx1678);
   ix20022 : mux21 port map ( Y=>nx20021, A0=>nx31914, A1=>nx42259, S0=>
      nx42271);
   ix31915 : aoi44 port map ( Y=>nx31914, A0=>nx42861, A1=>nx42259, A2=>
      nx41407, A3=>nx42865, B0=>nx31906, B1=>nx42877, B2=>nx41385, B3=>
      nx1602);
   ix18632 : mux21_ni port map ( Y=>nx18631, A0=>nx20, A1=>nx42861, S0=>
      nx42271);
   ix21 : oai21 port map ( Y=>nx20, A0=>nx42861, A1=>nx31919, B0=>nx31959);
   ix31920 : aoi21 port map ( Y=>nx31919, A0=>nx42259, A1=>nx42865, B0=>
      nx41377);
   ix20042 : nand02 port map ( Y=>nx20041, A0=>nx42877, A1=>nx42881);
   reg_state_2 : dffr port map ( Q=>state_2, QB=>OPEN, D=>nx20041, CLK=>clk, 
      R=>rst);
   ix1699 : nor03_2x port map ( Y=>nx18145, A0=>state_0, A1=>state_2, A2=>
      nx42883);
   reg_state_0 : dffr port map ( Q=>state_0, QB=>nx31906, D=>nx20051, CLK=>
      clk, R=>rst);
   ix20032 : oai22 port map ( Y=>nx20031, A0=>nx31933, A1=>nx32689, B0=>
      nx42883, B1=>nx42877);
   ix31934 : aoi221 port map ( Y=>nx31933, A0=>nx41391, A1=>nx18159, B0=>
      nx41375, B1=>nx31938, C0=>nx41389);
   reg_sub_state_2 : dffr port map ( Q=>sub_state_2, QB=>OPEN, D=>nx20021, 
      CLK=>clk, R=>rst);
   reg_state_1 : dffr port map ( Q=>OPEN, QB=>nx31930, D=>nx20031, CLK=>clk, 
      R=>rst);
   ix31939 : nand04 port map ( Y=>nx31938, A0=>nx742, A1=>nx1044, A2=>nx1348, 
      A3=>nx1576);
   ix743 : nor04 port map ( Y=>nx742, A0=>num_out_2, A1=>num_out_0, A2=>
      num_out_1, A3=>nx32202);
   num_loop1_2_fx_reg_q : dffr port map ( Q=>num_out_2, QB=>OPEN, D=>nx19101, 
      CLK=>clk, R=>rst);
   reg_num_in_2 : dff port map ( Q=>num_in_2, QB=>OPEN, D=>nx19091, CLK=>clk
   );
   ix31947 : xnor2 port map ( Y=>nx31946, A0=>nx31948, A1=>nx32175);
   ix31949 : aoi22 port map ( Y=>nx31948, A0=>nx41413, A1=>alu_inp1_1, B0=>
      nx442, B1=>nx18161);
   reg_alu_sel : dff port map ( Q=>alu_sel, QB=>OPEN, D=>nx18871, CLK=>clk);
   ix31956 : inv01 port map ( Y=>nx31955, A=>rst);
   ix31958 : aoi21 port map ( Y=>nx31957, A0=>nx31959, A1=>nx98, B0=>nx18155
   );
   ix31960 : nand02 port map ( Y=>nx31959, A0=>nx31961, A1=>nx41387);
   ix18642 : mux21_ni port map ( Y=>nx18641, A0=>nx50, A1=>nx41405, S0=>
      nx42271);
   ix51 : oai21 port map ( Y=>nx50, A0=>nx42249, A1=>nx31966, B0=>nx31968);
   ix31969 : oai21 port map ( Y=>nx31968, A0=>nx31970, A1=>nx31974, B0=>
      nx42865);
   reg_sub_state_1 : dffr port map ( Q=>OPEN, QB=>nx31972, D=>nx18641, CLK=>
      clk, R=>rst);
   reg_sub_state_0 : dffr port map ( Q=>sub_state_0, QB=>OPEN, D=>nx18631, 
      CLK=>clk, R=>rst);
   ix31979 : aoi21 port map ( Y=>nx31978, A0=>nx31938, A1=>nx1582, B0=>
      nx1592);
   ix18862 : nand02 port map ( Y=>nx18861, A0=>nx42897, A1=>nx43519);
   booth_shift_Reg_adder_0_reg_count_19 : dffr port map ( Q=>OPEN, QB=>
      nx31985, D=>nx18861, CLK=>clk, R=>nx42817);
   reg_ready_signal : dffr port map ( Q=>ready_signal, QB=>OPEN, D=>nx18661, 
      CLK=>clk, R=>rst);
   ix31992 : nand02 port map ( Y=>nx31991, A0=>nx31959, A1=>nx132);
   ix123 : nand03 port map ( Y=>nx122, A0=>nx42867, A1=>nx31961, A2=>nx31938
   );
   booth_shift_Reg_adder_0_reg_count_17 : dffr port map ( Q=>output_17, QB=>
      OPEN, D=>nx18841, CLK=>clk, R=>nx41473);
   booth_shift_Reg_adder_0_reg_count_16 : dffr port map ( Q=>output_16, QB=>
      OPEN, D=>nx18831, CLK=>clk, R=>nx41473);
   booth_shift_Reg_adder_0_reg_count_15 : dffr port map ( Q=>output_15, QB=>
      OPEN, D=>nx18821, CLK=>clk, R=>nx41473);
   booth_shift_Reg_adder_0_reg_count_14 : dffr port map ( Q=>output_14, QB=>
      OPEN, D=>nx18811, CLK=>clk, R=>nx41473);
   booth_shift_Reg_adder_0_reg_count_13 : dffr port map ( Q=>output_13, QB=>
      OPEN, D=>nx18801, CLK=>clk, R=>nx41473);
   booth_shift_Reg_adder_0_reg_count_12 : dffr port map ( Q=>output_12, QB=>
      OPEN, D=>nx18791, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_11 : dffr port map ( Q=>output_11, QB=>
      OPEN, D=>nx18781, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_10 : dffr port map ( Q=>output_10, QB=>
      OPEN, D=>nx18771, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_9 : dffr port map ( Q=>output_9, QB=>
      OPEN, D=>nx18761, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_8 : dffr port map ( Q=>output_8, QB=>
      OPEN, D=>nx18751, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_7 : dffr port map ( Q=>output_7, QB=>
      OPEN, D=>nx18741, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_6 : dffr port map ( Q=>output_6, QB=>
      OPEN, D=>nx18731, CLK=>clk, R=>nx41471);
   booth_shift_Reg_adder_0_reg_count_5 : dffr port map ( Q=>output_5, QB=>
      OPEN, D=>nx18721, CLK=>clk, R=>nx42817);
   booth_shift_Reg_adder_0_reg_count_4 : dffr port map ( Q=>output_4, QB=>
      OPEN, D=>nx18711, CLK=>clk, R=>nx42817);
   booth_shift_Reg_adder_0_reg_count_3 : dffr port map ( Q=>output_3, QB=>
      OPEN, D=>nx18701, CLK=>clk, R=>nx42817);
   booth_shift_Reg_adder_0_reg_count_2 : dffr port map ( Q=>output_2, QB=>
      OPEN, D=>nx18691, CLK=>clk, R=>nx42817);
   booth_shift_Reg_adder_0_reg_count_1 : dffr port map ( Q=>output_1, QB=>
      OPEN, D=>nx18681, CLK=>clk, R=>nx42817);
   booth_shift_Reg_adder_0_reg_count_0 : dffs_ni port map ( Q=>output_0, QB
      =>OPEN, D=>nx18667, CLK=>clk, S=>nx42817);
   ix18668 : nor02ii port map ( Y=>nx18667, A0=>nx42897, A1=>output_0);
   booth_shift_Reg_adder_0_reg_count_18 : dffr port map ( Q=>
      enable_decoder_dst_booth, QB=>OPEN, D=>nx18851, CLK=>clk, R=>nx41473);
   ix1593 : aoi21 port map ( Y=>nx1592, A0=>nx31906, A1=>nx41383, B0=>
      state_2);
   ix99 : nand02 port map ( Y=>nx98, A0=>nx18146, A1=>nx42277);
   ix247 : aoi22 port map ( Y=>nx246, A0=>nx42865, A1=>nx36, B0=>nx32062, B1
      =>nx41375);
   ix32063 : nand04 port map ( Y=>nx32062, A0=>nx42891, A1=>nx42867, A2=>
      nx42881, A3=>nx41405);
   reg_alu_inp1_1 : dff port map ( Q=>alu_inp1_1, QB=>OPEN, D=>nx19031, CLK
      =>clk);
   num_loop1_1_fx_reg_q : dffr port map ( Q=>num_out_1, QB=>OPEN, D=>nx19021, 
      CLK=>clk, R=>rst);
   ix32073 : aoi22 port map ( Y=>nx32072, A0=>data_in(1), A1=>nx41409, B0=>
      nx444, B1=>nx41387);
   ix445 : xnor2 port map ( Y=>nx444, A0=>nx442, A1=>nx32148);
   reg_alu_inp1_0 : dff port map ( Q=>alu_inp1_0, QB=>OPEN, D=>nx18951, CLK
      =>clk);
   num_loop1_0_fx_reg_q : dffr port map ( Q=>num_out_0, QB=>OPEN, D=>nx18941, 
      CLK=>clk, R=>rst);
   reg_num_in_0 : dff port map ( Q=>num_in_0, QB=>OPEN, D=>nx18931, CLK=>clk
   );
   reg_alu_inp2_0 : dff port map ( Q=>alu_inp2_0, QB=>nx32089, D=>nx18961, 
      CLK=>clk);
   ix18652 : nand02 port map ( Y=>nx18651, A0=>nx42907, A1=>nx32103);
   reg_enable_num : dffr port map ( Q=>OPEN, QB=>nx32101, D=>nx18651, CLK=>
      clk, R=>rst);
   ix32104 : nand02 port map ( Y=>nx32103, A0=>nx31961, A1=>nx41409);
   addr_loop1_0_fx_reg_q : dffr port map ( Q=>address_out(0), QB=>OPEN, D=>
      nx18921, CLK=>clk, R=>rst);
   reg_address_in_0 : dffr port map ( Q=>address_in_0, QB=>OPEN, D=>nx18911, 
      CLK=>clk, R=>rst);
   ix389 : oai22 port map ( Y=>nx388, A0=>nx32085, A1=>nx42313, B0=>nx42249, 
      B1=>nx32113);
   reg_neuron_address_0 : dffr port map ( Q=>neuron_address_0, QB=>OPEN, D=>
      nx18891, CLK=>clk, R=>rst);
   reg_temp_0 : dffr port map ( Q=>temp_0, QB=>OPEN, D=>nx18901, CLK=>clk, R
      =>rst);
   ix295 : aoi21 port map ( Y=>nx294, A0=>nx32119, A1=>nx18159, B0=>nx32126
   );
   ix32127 : aoi43 port map ( Y=>nx32126, A0=>nx41375, A1=>nx41391, A2=>
      nx42861, A3=>nx284, B0=>state_0, B1=>nx42877, B2=>nx42883);
   ix32132 : aoi332 port map ( Y=>nx32131, A0=>nx42299, A1=>nx42249, A2=>
      nx41515, B0=>nx338, B1=>nx42259, B2=>nx31966, C0=>nx306, C1=>nx326);
   ix339 : or02 port map ( Y=>nx338, A0=>nx336, A1=>nx41515);
   ix327 : aoi21 port map ( Y=>nx326, A0=>nx32119, A1=>nx18159, B0=>nx32137
   );
   ix32138 : aoi43 port map ( Y=>nx32137, A0=>nx42891, A1=>nx41375, A2=>
      nx42299, A3=>nx42887, B0=>nx31961, B1=>nx42877, B2=>nx42883);
   ix18882 : nand02 port map ( Y=>nx18881, A0=>nx42915, A1=>nx32144);
   reg_enable_address : dffr port map ( Q=>OPEN, QB=>nx32142, D=>nx18881, 
      CLK=>clk, R=>rst);
   ix32145 : nand02 port map ( Y=>nx32144, A0=>nx31974, A1=>nx41409);
   reg_num_in_1 : dff port map ( Q=>num_in_1, QB=>nx32150, D=>nx19011, CLK=>
      clk);
   addr_loop1_1_fx_reg_q : dffr port map ( Q=>address_out(1), QB=>OPEN, D=>
      nx19001, CLK=>clk, R=>rst);
   reg_address_in_1 : dffr port map ( Q=>address_in_1, QB=>OPEN, D=>nx18991, 
      CLK=>clk, R=>rst);
   ix18972 : oai21 port map ( Y=>nx18971, A0=>nx32164, A1=>nx41523, B0=>
      nx32166);
   reg_neuron_address_1 : dffr port map ( Q=>neuron_address_1, QB=>nx32164, 
      D=>nx18971, CLK=>clk, R=>rst);
   ix32167 : nand03 port map ( Y=>nx32166, A0=>nx41375, A1=>nx444, A2=>
      nx41523);
   reg_temp_1 : dffr port map ( Q=>temp_1, QB=>OPEN, D=>nx18981, CLK=>clk, R
      =>rst);
   reg_alu_inp1_2 : dff port map ( Q=>alu_inp1_2, QB=>nx32197, D=>nx19081, 
      CLK=>clk);
   addr_loop1_2_fx_reg_q : dffr port map ( Q=>address_out(2), QB=>OPEN, D=>
      nx19071, CLK=>clk, R=>rst);
   reg_address_in_2 : dffr port map ( Q=>address_in_2, QB=>OPEN, D=>nx19061, 
      CLK=>clk, R=>rst);
   ix539 : oai22 port map ( Y=>nx538, A0=>nx31946, A1=>nx42313, B0=>nx42251, 
      B1=>nx32185);
   reg_neuron_address_2 : dffr port map ( Q=>neuron_address_2, QB=>OPEN, D=>
      nx19041, CLK=>clk, R=>rst);
   reg_temp_2 : dffr port map ( Q=>temp_2, QB=>OPEN, D=>nx19051, CLK=>clk, R
      =>rst);
   ix32203 : or02 port map ( Y=>nx32202, A0=>num_out_3, A1=>num_out_4);
   num_loop1_3_fx_reg_q : dffr port map ( Q=>num_out_3, QB=>OPEN, D=>nx19171, 
      CLK=>clk, R=>rst);
   ix32209 : aoi22 port map ( Y=>nx32208, A0=>data_in(3), A1=>nx41409, B0=>
      nx18163, B1=>nx41387);
   ix647 : xnor2 port map ( Y=>nx18163, A0=>nx596, A1=>nx32212);
   ix597 : oai22 port map ( Y=>nx596, A0=>nx31948, A1=>nx32175, B0=>nx42295, 
      B1=>nx32197);
   reg_alu_inp1_3 : dff port map ( Q=>alu_inp1_3, QB=>OPEN, D=>nx19151, CLK
      =>clk);
   addr_loop1_3_fx_reg_q : dffr port map ( Q=>address_out(3), QB=>OPEN, D=>
      nx19141, CLK=>clk, R=>rst);
   reg_address_in_3 : dffr port map ( Q=>address_in_3, QB=>OPEN, D=>nx19131, 
      CLK=>clk, R=>rst);
   ix19112 : oai21 port map ( Y=>nx19111, A0=>nx32228, A1=>nx41523, B0=>
      nx32230);
   reg_neuron_address_3 : dffr port map ( Q=>neuron_address_3, QB=>nx32228, 
      D=>nx19111, CLK=>clk, R=>rst);
   ix32231 : nand03 port map ( Y=>nx32230, A0=>nx41375, A1=>nx18163, A2=>
      nx41523);
   reg_temp_3 : dffr port map ( Q=>temp_3, QB=>OPEN, D=>nx19121, CLK=>clk, R
      =>rst);
   reg_num_in_3 : dff port map ( Q=>num_in_3, QB=>nx32238, D=>nx19161, CLK=>
      clk);
   num_loop1_4_fx_reg_q : dffr port map ( Q=>num_out_4, QB=>OPEN, D=>nx19241, 
      CLK=>clk, R=>rst);
   reg_num_in_4 : dff port map ( Q=>num_in_4, QB=>OPEN, D=>nx19231, CLK=>clk
   );
   ix725 : oai22 port map ( Y=>nx724, A0=>nx32246, A1=>nx42279, B0=>nx32274, 
      B1=>nx42299);
   ix32247 : xnor2 port map ( Y=>nx32246, A0=>nx32248, A1=>nx32251);
   ix32249 : aoi22 port map ( Y=>nx32248, A0=>nx41413, A1=>alu_inp1_3, B0=>
      nx596, B1=>nx644);
   reg_alu_inp1_4 : dff port map ( Q=>alu_inp1_4, QB=>nx32273, D=>nx19221, 
      CLK=>clk);
   addr_loop1_4_fx_reg_q : dffr port map ( Q=>address_out(4), QB=>OPEN, D=>
      nx19211, CLK=>clk, R=>rst);
   reg_address_in_4 : dffr port map ( Q=>address_in_4, QB=>OPEN, D=>nx19201, 
      CLK=>clk, R=>rst);
   ix693 : oai22 port map ( Y=>nx692, A0=>nx32246, A1=>nx42313, B0=>nx42251, 
      B1=>nx32261);
   reg_neuron_address_4 : dffr port map ( Q=>neuron_address_4, QB=>OPEN, D=>
      nx19181, CLK=>clk, R=>rst);
   reg_temp_4 : dffr port map ( Q=>temp_4, QB=>OPEN, D=>nx19191, CLK=>clk, R
      =>rst);
   ix32275 : inv01 port map ( Y=>nx32274, A=>data_in(4));
   ix1045 : nor04 port map ( Y=>nx1044, A0=>num_out_5, A1=>num_out_6, A2=>
      num_out_7, A3=>num_out_8);
   num_loop1_5_fx_reg_q : dffr port map ( Q=>num_out_5, QB=>OPEN, D=>nx19311, 
      CLK=>clk, R=>rst);
   ix32284 : aoi22 port map ( Y=>nx32283, A0=>data_in(5), A1=>nx41411, B0=>
      nx18167, B1=>nx41387);
   ix799 : xnor2 port map ( Y=>nx18167, A0=>nx748, A1=>nx32287);
   ix749 : oai22 port map ( Y=>nx748, A0=>nx32248, A1=>nx32251, B0=>nx42295, 
      B1=>nx32273);
   reg_alu_inp1_5 : dff port map ( Q=>alu_inp1_5, QB=>OPEN, D=>nx19291, CLK
      =>clk);
   addr_loop1_5_fx_reg_q : dffr port map ( Q=>address_out(5), QB=>OPEN, D=>
      nx19281, CLK=>clk, R=>rst);
   reg_address_in_5 : dffr port map ( Q=>address_in_5, QB=>OPEN, D=>nx19271, 
      CLK=>clk, R=>rst);
   ix19252 : oai21 port map ( Y=>nx19251, A0=>nx32303, A1=>nx41525, B0=>
      nx32305);
   reg_neuron_address_5 : dffr port map ( Q=>neuron_address_5, QB=>nx32303, 
      D=>nx19251, CLK=>clk, R=>rst);
   ix32306 : nand03 port map ( Y=>nx32305, A0=>nx41377, A1=>nx18167, A2=>
      nx41525);
   reg_temp_5 : dffr port map ( Q=>temp_5, QB=>OPEN, D=>nx19261, CLK=>clk, R
      =>rst);
   reg_num_in_5 : dff port map ( Q=>num_in_5, QB=>nx32313, D=>nx19301, CLK=>
      clk);
   num_loop1_6_fx_reg_q : dffr port map ( Q=>num_out_6, QB=>OPEN, D=>nx19381, 
      CLK=>clk, R=>rst);
   reg_num_in_6 : dff port map ( Q=>num_in_6, QB=>OPEN, D=>nx19371, CLK=>clk
   );
   ix877 : oai22 port map ( Y=>nx876, A0=>nx32321, A1=>nx42279, B0=>nx32349, 
      B1=>nx42299);
   ix32322 : xnor2 port map ( Y=>nx32321, A0=>nx32323, A1=>nx32326);
   ix32324 : aoi22 port map ( Y=>nx32323, A0=>nx41415, A1=>alu_inp1_5, B0=>
      nx748, B1=>nx796);
   reg_alu_inp1_6 : dff port map ( Q=>alu_inp1_6, QB=>nx32348, D=>nx19361, 
      CLK=>clk);
   addr_loop1_6_fx_reg_q : dffr port map ( Q=>address_out(6), QB=>OPEN, D=>
      nx19351, CLK=>clk, R=>rst);
   reg_address_in_6 : dffr port map ( Q=>address_in_6, QB=>OPEN, D=>nx19341, 
      CLK=>clk, R=>rst);
   ix845 : oai22 port map ( Y=>nx844, A0=>nx32321, A1=>nx42313, B0=>nx42251, 
      B1=>nx32336);
   reg_neuron_address_6 : dffr port map ( Q=>neuron_address_6, QB=>OPEN, D=>
      nx19321, CLK=>clk, R=>rst);
   reg_temp_6 : dffr port map ( Q=>temp_6, QB=>OPEN, D=>nx19331, CLK=>clk, R
      =>rst);
   ix32350 : inv01 port map ( Y=>nx32349, A=>data_in(6));
   num_loop1_7_fx_reg_q : dffr port map ( Q=>num_out_7, QB=>OPEN, D=>nx19451, 
      CLK=>clk, R=>rst);
   ix32358 : aoi22 port map ( Y=>nx32357, A0=>data_in(7), A1=>nx41411, B0=>
      nx18171, B1=>nx41389);
   ix949 : xnor2 port map ( Y=>nx18171, A0=>nx898, A1=>nx32361);
   ix899 : oai22 port map ( Y=>nx898, A0=>nx32323, A1=>nx32326, B0=>nx42295, 
      B1=>nx32348);
   reg_alu_inp1_7 : dff port map ( Q=>alu_inp1_7, QB=>OPEN, D=>nx19431, CLK
      =>clk);
   addr_loop1_7_fx_reg_q : dffr port map ( Q=>address_out(7), QB=>OPEN, D=>
      nx19421, CLK=>clk, R=>rst);
   reg_address_in_7 : dffr port map ( Q=>address_in_7, QB=>OPEN, D=>nx19411, 
      CLK=>clk, R=>rst);
   ix19392 : oai21 port map ( Y=>nx19391, A0=>nx32377, A1=>nx41525, B0=>
      nx32379);
   reg_neuron_address_7 : dffr port map ( Q=>neuron_address_7, QB=>nx32377, 
      D=>nx19391, CLK=>clk, R=>rst);
   ix32380 : nand03 port map ( Y=>nx32379, A0=>nx41377, A1=>nx18171, A2=>
      nx41525);
   reg_temp_7 : dffr port map ( Q=>temp_7, QB=>OPEN, D=>nx19401, CLK=>clk, R
      =>rst);
   reg_num_in_7 : dff port map ( Q=>num_in_7, QB=>nx32387, D=>nx19441, CLK=>
      clk);
   num_loop1_8_fx_reg_q : dffr port map ( Q=>num_out_8, QB=>OPEN, D=>nx19521, 
      CLK=>clk, R=>rst);
   reg_num_in_8 : dff port map ( Q=>num_in_8, QB=>OPEN, D=>nx19511, CLK=>clk
   );
   ix1027 : oai22 port map ( Y=>nx1026, A0=>nx32395, A1=>nx42281, B0=>
      nx32423, B1=>nx42299);
   ix32396 : xnor2 port map ( Y=>nx32395, A0=>nx32397, A1=>nx32400);
   ix32398 : aoi22 port map ( Y=>nx32397, A0=>nx41415, A1=>alu_inp1_7, B0=>
      nx898, B1=>nx946);
   reg_alu_inp1_8 : dff port map ( Q=>alu_inp1_8, QB=>nx32422, D=>nx19501, 
      CLK=>clk);
   addr_loop1_8_fx_reg_q : dffr port map ( Q=>address_out(8), QB=>OPEN, D=>
      nx19491, CLK=>clk, R=>rst);
   reg_address_in_8 : dffr port map ( Q=>address_in_8, QB=>OPEN, D=>nx19481, 
      CLK=>clk, R=>rst);
   ix995 : oai22 port map ( Y=>nx994, A0=>nx32395, A1=>nx42315, B0=>nx42253, 
      B1=>nx32410);
   reg_neuron_address_8 : dffr port map ( Q=>neuron_address_8, QB=>OPEN, D=>
      nx19461, CLK=>clk, R=>rst);
   reg_temp_8 : dffr port map ( Q=>temp_8, QB=>OPEN, D=>nx19471, CLK=>clk, R
      =>rst);
   ix32424 : inv01 port map ( Y=>nx32423, A=>data_in(8));
   ix1349 : nor04 port map ( Y=>nx1348, A0=>num_out_9, A1=>num_out_10, A2=>
      num_out_11, A3=>num_out_12);
   num_loop1_9_fx_reg_q : dffr port map ( Q=>num_out_9, QB=>OPEN, D=>nx19591, 
      CLK=>clk, R=>rst);
   ix32433 : aoi22 port map ( Y=>nx32432, A0=>data_in(9), A1=>nx41411, B0=>
      nx18175, B1=>nx41389);
   ix1103 : xnor2 port map ( Y=>nx18175, A0=>nx1052, A1=>nx32436);
   ix1053 : oai22 port map ( Y=>nx1052, A0=>nx32397, A1=>nx32400, B0=>
      nx42295, B1=>nx32422);
   reg_alu_inp1_9 : dff port map ( Q=>alu_inp1_9, QB=>OPEN, D=>nx19571, CLK
      =>clk);
   addr_loop1_9_fx_reg_q : dffr port map ( Q=>address_out(9), QB=>OPEN, D=>
      nx19561, CLK=>clk, R=>rst);
   reg_address_in_9 : dffr port map ( Q=>address_in_9, QB=>OPEN, D=>nx19551, 
      CLK=>clk, R=>rst);
   ix19532 : oai21 port map ( Y=>nx19531, A0=>nx32452, A1=>nx41525, B0=>
      nx32454);
   reg_neuron_address_9 : dffr port map ( Q=>neuron_address_9, QB=>nx32452, 
      D=>nx19531, CLK=>clk, R=>rst);
   ix32455 : nand03 port map ( Y=>nx32454, A0=>nx41377, A1=>nx18175, A2=>
      nx41527);
   reg_temp_9 : dffr port map ( Q=>temp_9, QB=>OPEN, D=>nx19541, CLK=>clk, R
      =>rst);
   reg_num_in_9 : dff port map ( Q=>num_in_9, QB=>nx32462, D=>nx19581, CLK=>
      clk);
   num_loop1_10_fx_reg_q : dffr port map ( Q=>num_out_10, QB=>OPEN, D=>
      nx19661, CLK=>clk, R=>rst);
   reg_num_in_10 : dff port map ( Q=>num_in_10, QB=>OPEN, D=>nx19651, CLK=>
      clk);
   ix1181 : oai22 port map ( Y=>nx1180, A0=>nx32470, A1=>nx42281, B0=>
      nx32498, B1=>nx43103);
   ix32471 : xnor2 port map ( Y=>nx32470, A0=>nx32472, A1=>nx32475);
   ix32473 : aoi22 port map ( Y=>nx32472, A0=>nx41417, A1=>alu_inp1_9, B0=>
      nx1052, B1=>nx1100);
   reg_alu_inp1_10 : dff port map ( Q=>alu_inp1_10, QB=>nx32497, D=>nx19641, 
      CLK=>clk);
   addr_loop1_10_fx_reg_q : dffr port map ( Q=>address_out(10), QB=>OPEN, D
      =>nx19631, CLK=>clk, R=>rst);
   reg_address_in_10 : dffr port map ( Q=>address_in_10, QB=>OPEN, D=>
      nx19621, CLK=>clk, R=>rst);
   ix1149 : oai22 port map ( Y=>nx1148, A0=>nx32470, A1=>nx42315, B0=>
      nx42253, B1=>nx32485);
   reg_neuron_address_10 : dffr port map ( Q=>neuron_address_10, QB=>OPEN, D
      =>nx19601, CLK=>clk, R=>rst);
   reg_temp_10 : dffr port map ( Q=>temp_10, QB=>OPEN, D=>nx19611, CLK=>clk, 
      R=>rst);
   ix32499 : inv01 port map ( Y=>nx32498, A=>data_in(10));
   num_loop1_11_fx_reg_q : dffr port map ( Q=>num_out_11, QB=>OPEN, D=>
      nx19731, CLK=>clk, R=>rst);
   ix32507 : aoi22 port map ( Y=>nx32506, A0=>data_in(11), A1=>nx41411, B0=>
      nx18178, B1=>nx41389);
   ix1253 : xnor2 port map ( Y=>nx18178, A0=>nx1202, A1=>nx32510);
   ix1203 : oai22 port map ( Y=>nx1202, A0=>nx32472, A1=>nx32475, B0=>
      nx42295, B1=>nx32497);
   reg_alu_inp1_11 : dff port map ( Q=>alu_inp1_11, QB=>OPEN, D=>nx19711, 
      CLK=>clk);
   addr_loop1_11_fx_reg_q : dffr port map ( Q=>address_out(11), QB=>OPEN, D
      =>nx19701, CLK=>clk, R=>rst);
   reg_address_in_11 : dffr port map ( Q=>address_in_11, QB=>OPEN, D=>
      nx19691, CLK=>clk, R=>rst);
   ix19672 : oai21 port map ( Y=>nx19671, A0=>nx32526, A1=>nx41527, B0=>
      nx32528);
   reg_neuron_address_11 : dffr port map ( Q=>neuron_address_11, QB=>nx32526, 
      D=>nx19671, CLK=>clk, R=>rst);
   ix32529 : nand03 port map ( Y=>nx32528, A0=>nx41377, A1=>nx18178, A2=>
      nx41527);
   reg_temp_11 : dffr port map ( Q=>temp_11, QB=>OPEN, D=>nx19681, CLK=>clk, 
      R=>rst);
   reg_num_in_11 : dff port map ( Q=>num_in_11, QB=>nx32536, D=>nx19721, CLK
      =>clk);
   num_loop1_12_fx_reg_q : dffr port map ( Q=>num_out_12, QB=>OPEN, D=>
      nx19801, CLK=>clk, R=>rst);
   reg_num_in_12 : dff port map ( Q=>num_in_12, QB=>OPEN, D=>nx19791, CLK=>
      clk);
   ix1331 : oai22 port map ( Y=>nx1330, A0=>nx32544, A1=>nx42283, B0=>
      nx32572, B1=>nx43103);
   ix32545 : xnor2 port map ( Y=>nx32544, A0=>nx32546, A1=>nx32549);
   ix32547 : aoi22 port map ( Y=>nx32546, A0=>nx41417, A1=>alu_inp1_11, B0=>
      nx1202, B1=>nx1250);
   reg_alu_inp1_12 : dff port map ( Q=>alu_inp1_12, QB=>nx32571, D=>nx19781, 
      CLK=>clk);
   addr_loop1_12_fx_reg_q : dffr port map ( Q=>address_out(12), QB=>OPEN, D
      =>nx19771, CLK=>clk, R=>rst);
   reg_address_in_12 : dffr port map ( Q=>address_in_12, QB=>OPEN, D=>
      nx19761, CLK=>clk, R=>rst);
   ix1299 : oai22 port map ( Y=>nx1298, A0=>nx32544, A1=>nx42315, B0=>
      nx42255, B1=>nx32559);
   reg_neuron_address_12 : dffr port map ( Q=>neuron_address_12, QB=>OPEN, D
      =>nx19741, CLK=>clk, R=>rst);
   reg_temp_12 : dffr port map ( Q=>temp_12, QB=>OPEN, D=>nx19751, CLK=>clk, 
      R=>rst);
   ix32573 : inv01 port map ( Y=>nx32572, A=>data_in(12));
   ix1577 : nor04 port map ( Y=>nx1576, A0=>num_out_13, A1=>num_out_14, A2=>
      num_out_15, A3=>nx42897);
   num_loop1_13_fx_reg_q : dffr port map ( Q=>num_out_13, QB=>OPEN, D=>
      nx19871, CLK=>clk, R=>rst);
   ix32582 : aoi22 port map ( Y=>nx32581, A0=>data_in(13), A1=>nx41411, B0=>
      nx18180, B1=>nx41389);
   ix1405 : xnor2 port map ( Y=>nx18180, A0=>nx1354, A1=>nx32585);
   ix1355 : oai22 port map ( Y=>nx1354, A0=>nx32546, A1=>nx32549, B0=>
      nx42295, B1=>nx32571);
   reg_alu_inp1_13 : dff port map ( Q=>alu_inp1_13, QB=>OPEN, D=>nx19851, 
      CLK=>clk);
   addr_loop1_13_fx_reg_q : dffr port map ( Q=>address_out(13), QB=>OPEN, D
      =>nx19841, CLK=>clk, R=>rst);
   reg_address_in_13 : dffr port map ( Q=>address_in_13, QB=>OPEN, D=>
      nx19831, CLK=>clk, R=>rst);
   ix19812 : oai21 port map ( Y=>nx19811, A0=>nx32601, A1=>nx41527, B0=>
      nx32603);
   reg_neuron_address_13 : dffr port map ( Q=>neuron_address_13, QB=>nx32601, 
      D=>nx19811, CLK=>clk, R=>rst);
   ix32604 : nand03 port map ( Y=>nx32603, A0=>nx41377, A1=>nx18180, A2=>
      nx41527);
   reg_temp_13 : dffr port map ( Q=>temp_13, QB=>OPEN, D=>nx19821, CLK=>clk, 
      R=>rst);
   reg_num_in_13 : dff port map ( Q=>num_in_13, QB=>nx32611, D=>nx19861, CLK
      =>clk);
   num_loop1_14_fx_reg_q : dffr port map ( Q=>num_out_14, QB=>OPEN, D=>
      nx19941, CLK=>clk, R=>rst);
   reg_num_in_14 : dff port map ( Q=>num_in_14, QB=>OPEN, D=>nx19931, CLK=>
      clk);
   ix1483 : oai22 port map ( Y=>nx1482, A0=>nx32619, A1=>nx42283, B0=>
      nx32647, B1=>nx43103);
   ix32620 : xnor2 port map ( Y=>nx32619, A0=>nx32621, A1=>nx32624);
   ix32622 : aoi22 port map ( Y=>nx32621, A0=>nx41419, A1=>alu_inp1_13, B0=>
      nx1354, B1=>nx1402);
   reg_alu_inp1_14 : dff port map ( Q=>alu_inp1_14, QB=>nx32646, D=>nx19921, 
      CLK=>clk);
   addr_loop1_14_fx_reg_q : dffr port map ( Q=>address_out(14), QB=>OPEN, D
      =>nx19911, CLK=>clk, R=>rst);
   reg_address_in_14 : dffr port map ( Q=>address_in_14, QB=>OPEN, D=>
      nx19901, CLK=>clk, R=>rst);
   ix1451 : oai22 port map ( Y=>nx1450, A0=>nx32619, A1=>nx42317, B0=>
      nx42255, B1=>nx32634);
   reg_neuron_address_14 : dffr port map ( Q=>neuron_address_14, QB=>OPEN, D
      =>nx19881, CLK=>clk, R=>rst);
   reg_temp_14 : dffr port map ( Q=>temp_14, QB=>OPEN, D=>nx19891, CLK=>clk, 
      R=>rst);
   ix32648 : inv01 port map ( Y=>nx32647, A=>data_in(14));
   num_loop1_15_fx_reg_q : dffr port map ( Q=>num_out_15, QB=>OPEN, D=>
      nx20011, CLK=>clk, R=>rst);
   ix32656 : aoi22 port map ( Y=>nx32655, A0=>data_in(15), A1=>nx41411, B0=>
      nx18182, B1=>nx41389);
   ix1555 : xnor2 port map ( Y=>nx18182, A0=>nx1504, A1=>nx32659);
   ix1505 : oai22 port map ( Y=>nx1504, A0=>nx32621, A1=>nx32624, B0=>
      nx42295, B1=>nx32646);
   reg_alu_inp1_15 : dff port map ( Q=>alu_inp1_15, QB=>OPEN, D=>nx19991, 
      CLK=>clk);
   addr_loop1_15_fx_reg_q : dffr port map ( Q=>address_out(15), QB=>OPEN, D
      =>nx19981, CLK=>clk, R=>rst);
   reg_address_in_15 : dffr port map ( Q=>address_in_15, QB=>OPEN, D=>
      nx19971, CLK=>clk, R=>rst);
   ix19952 : oai21 port map ( Y=>nx19951, A0=>nx32676, A1=>nx41529, B0=>
      nx32678);
   reg_neuron_address_15 : dffr port map ( Q=>neuron_address_15, QB=>nx32676, 
      D=>nx19951, CLK=>clk, R=>rst);
   ix32679 : nand03 port map ( Y=>nx32678, A0=>nx18182, A1=>nx41377, A2=>
      nx41529);
   reg_temp_15 : dffr port map ( Q=>temp_15, QB=>OPEN, D=>nx19961, CLK=>clk, 
      R=>rst);
   reg_num_in_15 : dff port map ( Q=>num_in_15, QB=>nx32686, D=>nx20001, CLK
      =>clk);
   ix1603 : nand02 port map ( Y=>nx1602, A0=>nx32693, A1=>nx32119);
   ix32694 : oai21 port map ( Y=>nx32693, A0=>nx42891, A1=>nx42887, B0=>
      nx41397);
   ix1679 : aoi21 port map ( Y=>nx1678, A0=>nx32696, A1=>nx43103, B0=>
      nx43041);
   ix32697 : nand04 port map ( Y=>nx32696, A0=>nx41379, A1=>nx41407, A2=>
      nx42861, A3=>nx1672);
   ix32701 : aoi32 port map ( Y=>nx32700, A0=>max_calc_state_0, A1=>nx41563, 
      A2=>nx41313, B0=>nx33447, B1=>nx41585);
   ix20092 : mux21_ni port map ( Y=>nx20091, A0=>nx1774, A1=>
      max_calc_state_0, S0=>nx33444);
   ix1775 : nand03 port map ( Y=>nx1774, A0=>nx32705, A1=>nx31899, A2=>
      nx41310);
   ix32710 : nor02ii port map ( Y=>nx32709, A0=>nx32711, A1=>nx41031);
   ix32712 : nor04 port map ( Y=>nx32711, A0=>nx20306, A1=>nx20292, A2=>
      nx20276, A3=>nx20262);
   ix20307 : nand04 port map ( Y=>nx20306, A0=>nx32714, A1=>nx40998, A2=>
      nx41000, A3=>nx41002);
   max_calc_reg_answer_15 : dffr port map ( Q=>max_calc_answer_15, QB=>OPEN, 
      D=>nx31811, CLK=>clk, R=>rst);
   max_calc_reg_comparator_first_inp1_15 : dff port map ( Q=>
      max_calc_comparator_first_inp1_15, QB=>OPEN, D=>nx31621, CLK=>clk);
   lat_label_1_input_15 : latch port map ( Q=>label_1_input_15, D=>nx20006, 
      CLK=>nx41665);
   reg_label_1_input_state_machine_15 : dffr port map ( Q=>
      label_1_input_state_machine_15, QB=>OPEN, D=>nx31571, CLK=>clk, R=>rst
   );
   ix32730 : nand02 port map ( Y=>nx32729, A0=>nx41397, A1=>nx18159);
   ix20003 : xnor2 port map ( Y=>nx20002, A0=>nx32733, A1=>nx20000);
   ix32734 : aoi22 port map ( Y=>nx32733, A0=>label_1_output_14, A1=>
      booth_booth_integration_output_0_26, B0=>nx18050, B1=>nx18052);
   labelsregfile_label1_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_1_output_14, QB=>OPEN, D=>nx30381, CLK=>clk, R=>rst);
   lat_label_1_input_14 : latch port map ( Q=>label_1_input_14, D=>nx18058, 
      CLK=>nx41665);
   reg_label_1_input_state_machine_14 : dffr port map ( Q=>
      label_1_input_state_machine_14, QB=>OPEN, D=>nx30111, CLK=>clk, R=>rst
   );
   ix18055 : xnor2 port map ( Y=>nx18054, A0=>nx18050, A1=>nx33416);
   ix18051 : oai22 port map ( Y=>nx18050, A0=>nx32744, A1=>nx33405, B0=>
      nx33415, B1=>nx33152);
   ix32745 : aoi22 port map ( Y=>nx32744, A0=>label_1_output_12, A1=>
      booth_booth_integration_output_0_24, B0=>nx17986, B1=>nx18599);
   labelsregfile_label1_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_1_output_12, QB=>OPEN, D=>nx30351, CLK=>clk, R=>rst);
   lat_label_1_input_12 : latch port map ( Q=>label_1_input_12, D=>nx18000, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_12 : dffr port map ( Q=>
      label_1_input_state_machine_12, QB=>OPEN, D=>nx30341, CLK=>clk, R=>rst
   );
   ix17997 : xnor2 port map ( Y=>nx17996, A0=>nx17986, A1=>nx33401);
   ix17987 : oai22 port map ( Y=>nx17986, A0=>nx32755, A1=>nx33390, B0=>
      nx33400, B1=>nx33118);
   ix32756 : aoi22 port map ( Y=>nx32755, A0=>label_1_output_10, A1=>
      booth_booth_integration_output_0_22, B0=>nx17922, B1=>nx18597);
   labelsregfile_label1_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_1_output_10, QB=>OPEN, D=>nx30311, CLK=>clk, R=>rst);
   lat_label_1_input_10 : latch port map ( Q=>label_1_input_10, D=>nx17936, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_10 : dffr port map ( Q=>
      label_1_input_state_machine_10, QB=>OPEN, D=>nx30301, CLK=>clk, R=>rst
   );
   ix17933 : xnor2 port map ( Y=>nx17932, A0=>nx17922, A1=>nx33386);
   ix17923 : oai22 port map ( Y=>nx17922, A0=>nx32766, A1=>nx33375, B0=>
      nx33385, B1=>nx33084);
   ix32767 : aoi22 port map ( Y=>nx32766, A0=>label_1_output_8, A1=>
      booth_booth_integration_output_0_20, B0=>nx17858, B1=>nx18595);
   labelsregfile_label1_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_1_output_8, QB=>OPEN, D=>nx30271, CLK=>clk, R=>rst);
   lat_label_1_input_8 : latch port map ( Q=>label_1_input_8, D=>nx17872, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_8 : dffr port map ( Q=>
      label_1_input_state_machine_8, QB=>OPEN, D=>nx30261, CLK=>clk, R=>rst
   );
   ix17869 : xnor2 port map ( Y=>nx17868, A0=>nx17858, A1=>nx33371);
   ix17859 : oai22 port map ( Y=>nx17858, A0=>nx32777, A1=>nx33360, B0=>
      nx33370, B1=>nx33048);
   ix32778 : aoi22 port map ( Y=>nx32777, A0=>label_1_output_6, A1=>
      booth_booth_integration_output_0_18, B0=>nx17794, B1=>nx18593);
   labelsregfile_label1_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_1_output_6, QB=>OPEN, D=>nx30231, CLK=>clk, R=>rst);
   lat_label_1_input_6 : latch port map ( Q=>label_1_input_6, D=>nx17808, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_6 : dffr port map ( Q=>
      label_1_input_state_machine_6, QB=>OPEN, D=>nx30221, CLK=>clk, R=>rst
   );
   ix17805 : xnor2 port map ( Y=>nx17804, A0=>nx17794, A1=>nx33356);
   ix17795 : oai22 port map ( Y=>nx17794, A0=>nx32788, A1=>nx33345, B0=>
      nx33355, B1=>nx33011);
   ix32789 : aoi22 port map ( Y=>nx32788, A0=>label_1_output_4, A1=>
      booth_booth_integration_output_0_16, B0=>nx17730, B1=>nx18589);
   labelsregfile_label1_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_1_output_4, QB=>OPEN, D=>nx30191, CLK=>clk, R=>rst);
   lat_label_1_input_4 : latch port map ( Q=>label_1_input_4, D=>nx17744, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_4 : dffr port map ( Q=>
      label_1_input_state_machine_4, QB=>OPEN, D=>nx30181, CLK=>clk, R=>rst
   );
   ix17741 : xnor2 port map ( Y=>nx17740, A0=>nx17730, A1=>nx33341);
   ix17731 : oai22 port map ( Y=>nx17730, A0=>nx32799, A1=>nx33330, B0=>
      nx33340, B1=>nx33280);
   ix32800 : aoi22 port map ( Y=>nx32799, A0=>label_1_output_2, A1=>
      booth_booth_integration_output_0_14, B0=>nx17666, B1=>nx18585);
   labelsregfile_label1_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_1_output_2, QB=>OPEN, D=>nx30151, CLK=>clk, R=>rst);
   lat_label_1_input_2 : latch port map ( Q=>label_1_input_2, D=>nx17680, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_2 : dffr port map ( Q=>
      label_1_input_state_machine_2, QB=>OPEN, D=>nx30141, CLK=>clk, R=>rst
   );
   ix17677 : xnor2 port map ( Y=>nx17676, A0=>nx17666, A1=>nx33326);
   ix17667 : oai22 port map ( Y=>nx17666, A0=>nx32810, A1=>nx33315, B0=>
      nx33325, B1=>nx33289);
   ix32811 : nand02 port map ( Y=>nx32810, A0=>label_1_output_0, A1=>
      booth_booth_integration_output_0_12);
   labelsregfile_label1_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_1_output_0, QB=>OPEN, D=>nx20821, CLK=>clk, R=>rst);
   lat_label_1_input_0 : latch port map ( Q=>label_1_input_0, D=>nx2830, CLK
      =>nx41661);
   ix2831 : oai21 port map ( Y=>nx2830, A0=>nx32816, A1=>nx41421, B0=>
      nx32820);
   reg_label_1_input_state_machine_0 : dffr port map ( Q=>
      label_1_input_state_machine_0, QB=>nx32816, D=>nx20811, CLK=>clk, R=>
      rst);
   ix32821 : oai21 port map ( Y=>nx32820, A0=>
      booth_booth_integration_output_0_12, A1=>label_1_output_0, B0=>nx2818
   );
   booth_booth_integrtaion_0_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_12, QB=>OPEN, D=>nx20801, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_13, QB=>nx33289, D=>nx20781, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_14, QB=>OPEN, D=>nx20761, CLK=>clk, R
      =>rst);
   ix32834 : aoi22 port map ( Y=>nx32833, A0=>nx41795, A1=>nx41721, B0=>
      nx2734, B1=>nx2740);
   reg_neuron_15 : dff port map ( Q=>neuron_15, QB=>OPEN, D=>nx20731, CLK=>
      clk);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_reg_output_0, QB=>OPEN, 
      D=>nx20141, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_0, QB=>OPEN, D=>nx20127, CLK
      =>clk, S=>nx41477);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_reg_output_9, QB=>OPEN, 
      D=>nx20321, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_9, QB=>OPEN, D=>nx20311, CLK
      =>clk, R=>nx41477);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12688, QB=>OPEN, D=>nx20301, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_8, QB=>OPEN, D=>nx20291, CLK
      =>clk, R=>nx41477);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12689, QB=>OPEN, D=>nx20281, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_7, QB=>OPEN, D=>nx20271, CLK
      =>clk, R=>nx41477);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12690, QB=>OPEN, D=>nx20261, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_6, QB=>OPEN, D=>nx20251, CLK
      =>clk, R=>nx41475);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12691, QB=>OPEN, D=>nx20241, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_5, QB=>OPEN, D=>nx20231, CLK
      =>clk, R=>nx41475);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12692, QB=>OPEN, D=>nx20221, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_4, QB=>OPEN, D=>nx20211, CLK
      =>clk, R=>nx41475);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12693, QB=>OPEN, D=>nx20201, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_3, QB=>OPEN, D=>nx20191, CLK
      =>clk, R=>nx41475);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12694, QB=>OPEN, D=>nx20181, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_2, QB=>OPEN, D=>nx20171, CLK
      =>clk, R=>nx41475);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12695, QB=>OPEN, D=>nx20161, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_1, QB=>OPEN, D=>nx20151, CLK
      =>clk, R=>nx41475);
   ix20122 : nand02 port map ( Y=>nx20121, A0=>nx42921, A1=>nx41707);
   booth_booth_integrtaion_0_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx32886, D=>nx20121, CLK=>clk, S=>nx41475);
   ix2735 : nand02 port map ( Y=>nx2734, A0=>nx32907, A1=>nx33001);
   ix32908 : oai21 port map ( Y=>nx32907, A0=>nx41789, A1=>nx41785, B0=>
      data_in(0));
   ix20572 : oai21 port map ( Y=>nx20571, A0=>nx32912, A1=>nx42373, B0=>
      nx32914);
   booth_booth_integrtaion_0_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx32912, D=>nx20571, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0, QB=>nx32999, D=>nx20561, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1, QB=>OPEN, D=>nx20541, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2, QB=>OPEN, D=>nx20521, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3, QB=>OPEN, D=>nx20501, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4, QB=>OPEN, D=>nx20481, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5, QB=>OPEN, D=>nx20461, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6, QB=>OPEN, D=>nx20441, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7, QB=>OPEN, D=>nx20421, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8, QB=>OPEN, D=>nx20401, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9, QB=>OPEN, D=>nx20381, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10, QB=>OPEN, D=>nx20361, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11, QB=>OPEN, D=>nx20341, CLK=>clk, R=>rst);
   reg_neuron_11 : dff port map ( Q=>neuron_11, QB=>OPEN, D=>nx20331, CLK=>
      clk);
   reg_neuron_10 : dff port map ( Q=>neuron_10, QB=>OPEN, D=>nx20351, CLK=>
      clk);
   reg_neuron_9 : dff port map ( Q=>neuron_9, QB=>OPEN, D=>nx20371, CLK=>clk
   );
   reg_neuron_8 : dff port map ( Q=>neuron_8, QB=>OPEN, D=>nx20391, CLK=>clk
   );
   reg_neuron_7 : dff port map ( Q=>neuron_7, QB=>OPEN, D=>nx20411, CLK=>clk
   );
   reg_neuron_6 : dff port map ( Q=>neuron_6, QB=>OPEN, D=>nx20431, CLK=>clk
   );
   reg_neuron_5 : dff port map ( Q=>neuron_5, QB=>OPEN, D=>nx20451, CLK=>clk
   );
   reg_neuron_4 : dff port map ( Q=>neuron_4, QB=>OPEN, D=>nx20471, CLK=>clk
   );
   reg_neuron_3 : dff port map ( Q=>neuron_3, QB=>OPEN, D=>nx20491, CLK=>clk
   );
   reg_neuron_2 : dff port map ( Q=>neuron_2, QB=>OPEN, D=>nx20511, CLK=>clk
   );
   reg_neuron_1 : dff port map ( Q=>neuron_1, QB=>OPEN, D=>nx20531, CLK=>clk
   );
   reg_neuron_0 : dff port map ( Q=>neuron_0, QB=>OPEN, D=>nx20551, CLK=>clk
   );
   ix33006 : xnor2 port map ( Y=>nx33005, A0=>nx2204, A1=>nx18195);
   ix20712 : oai21 port map ( Y=>nx20711, A0=>nx33011, A1=>nx42373, B0=>
      nx33013);
   booth_booth_integrtaion_0_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_17, QB=>nx33011, D=>nx20711, CLK=>clk, 
      R=>rst);
   ix33014 : nand03 port map ( Y=>nx33013, A0=>nx42381, A1=>nx2712, A2=>
      nx42377);
   ix2713 : xnor2 port map ( Y=>nx2712, A0=>nx33016, A1=>nx18196);
   ix33017 : aoi22 port map ( Y=>nx33016, A0=>
      booth_booth_integration_output_0_17, A1=>nx2228, B0=>nx2204, B1=>
      nx18195);
   ix2219 : nor02_2x port map ( Y=>nx2218, A0=>data_in(0), A1=>data_in(1));
   ix20702 : oai21 port map ( Y=>nx20701, A0=>nx33031, A1=>nx42373, B0=>
      nx33033);
   booth_booth_integrtaion_0_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_18, QB=>nx33031, D=>nx20701, CLK=>clk, 
      R=>rst);
   ix33034 : nand03 port map ( Y=>nx33033, A0=>nx42381, A1=>nx2700, A2=>
      nx42377);
   ix2701 : xnor2 port map ( Y=>nx2700, A0=>nx2256, A1=>nx33044);
   ix2257 : oai22 port map ( Y=>nx2256, A0=>nx33016, A1=>nx33037, B0=>
      nx33031, B1=>nx42385);
   ix33040 : aoi32 port map ( Y=>nx33039, A0=>nx2238, A1=>nx41789, A2=>
      nx33042, B0=>data_in(2), B1=>nx41785);
   ix2239 : oai21 port map ( Y=>nx2238, A0=>data_in(0), A1=>data_in(1), B0=>
      data_in(2));
   ix20692 : oai21 port map ( Y=>nx20691, A0=>nx33048, A1=>nx42373, B0=>
      nx33050);
   booth_booth_integrtaion_0_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_19, QB=>nx33048, D=>nx20691, CLK=>clk, 
      R=>rst);
   ix33051 : nand03 port map ( Y=>nx33050, A0=>nx42381, A1=>nx2688, A2=>
      nx42377);
   ix2689 : xnor2 port map ( Y=>nx2688, A0=>nx33053, A1=>nx18198);
   ix33054 : aoi22 port map ( Y=>nx33053, A0=>
      booth_booth_integration_output_0_19, A1=>nx2276, B0=>nx2256, B1=>
      nx18197);
   ix2277 : oai32 port map ( Y=>nx2276, A0=>nx33056, A1=>nx33023, A2=>nx2266, 
      B0=>nx33059, B1=>nx33026);
   ix2243 : nor03_2x port map ( Y=>nx2242, A0=>data_in(2), A1=>data_in(0), 
      A2=>data_in(1));
   ix33060 : inv01 port map ( Y=>nx33059, A=>data_in(3));
   ix2267 : nor04 port map ( Y=>nx2266, A0=>data_in(3), A1=>data_in(2), A2=>
      data_in(0), A3=>data_in(1));
   ix33068 : xnor2 port map ( Y=>nx33067, A0=>nx2304, A1=>nx18199);
   ix2305 : oai22 port map ( Y=>nx2304, A0=>nx33053, A1=>nx33070, B0=>
      nx33079, B1=>nx42387);
   ix33073 : aoi32 port map ( Y=>nx33072, A0=>nx2286, A1=>nx41789, A2=>
      nx33077, B0=>data_in(4), B1=>nx41785);
   ix2287 : nand02 port map ( Y=>nx2286, A0=>nx33075, A1=>data_in(4));
   ix33078 : nand02 port map ( Y=>nx33077, A0=>nx32274, A1=>nx2266);
   booth_booth_integrtaion_0_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_20, QB=>nx33079, D=>nx20681, CLK=>clk, 
      R=>rst);
   ix20672 : oai21 port map ( Y=>nx20671, A0=>nx33084, A1=>nx42373, B0=>
      nx33086);
   booth_booth_integrtaion_0_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_21, QB=>nx33084, D=>nx20671, CLK=>clk, 
      R=>rst);
   ix33087 : nand03 port map ( Y=>nx33086, A0=>nx42381, A1=>nx2664, A2=>
      nx42377);
   ix2665 : xnor2 port map ( Y=>nx2664, A0=>nx33089, A1=>nx18200);
   ix33090 : aoi22 port map ( Y=>nx33089, A0=>
      booth_booth_integration_output_0_21, A1=>nx2324, B0=>nx2304, B1=>
      nx18199);
   ix2315 : nor02_2x port map ( Y=>nx2314, A0=>data_in(5), A1=>nx33077);
   ix33102 : xnor2 port map ( Y=>nx33101, A0=>nx2352, A1=>nx18201);
   ix2353 : oai22 port map ( Y=>nx2352, A0=>nx33089, A1=>nx33104, B0=>
      nx33113, B1=>nx42389);
   ix33107 : aoi32 port map ( Y=>nx33106, A0=>nx2334, A1=>nx41789, A2=>
      nx33111, B0=>data_in(6), B1=>nx41785);
   ix2335 : nand02 port map ( Y=>nx2334, A0=>nx33109, A1=>data_in(6));
   ix33112 : nand02 port map ( Y=>nx33111, A0=>nx32349, A1=>nx2314);
   booth_booth_integrtaion_0_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_22, QB=>nx33113, D=>nx20661, CLK=>clk, 
      R=>rst);
   ix20652 : oai21 port map ( Y=>nx20651, A0=>nx33118, A1=>nx42375, B0=>
      nx33120);
   booth_booth_integrtaion_0_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_23, QB=>nx33118, D=>nx20651, CLK=>clk, 
      R=>rst);
   ix33121 : nand03 port map ( Y=>nx33120, A0=>nx42381, A1=>nx2640, A2=>
      nx42377);
   ix2641 : xnor2 port map ( Y=>nx2640, A0=>nx33123, A1=>nx18203);
   ix33124 : aoi22 port map ( Y=>nx33123, A0=>
      booth_booth_integration_output_0_23, A1=>nx2372, B0=>nx2352, B1=>
      nx18201);
   ix2363 : nor02_2x port map ( Y=>nx2362, A0=>data_in(7), A1=>nx33111);
   ix33136 : xnor2 port map ( Y=>nx33135, A0=>nx2400, A1=>nx18205);
   ix2401 : oai22 port map ( Y=>nx2400, A0=>nx33123, A1=>nx33138, B0=>
      nx33147, B1=>nx42391);
   ix33141 : aoi32 port map ( Y=>nx33140, A0=>nx2382, A1=>nx41789, A2=>
      nx33145, B0=>data_in(8), B1=>nx41785);
   ix2383 : nand02 port map ( Y=>nx2382, A0=>nx33143, A1=>data_in(8));
   ix33146 : nand02 port map ( Y=>nx33145, A0=>nx32423, A1=>nx2362);
   booth_booth_integrtaion_0_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_24, QB=>nx33147, D=>nx20641, CLK=>clk, 
      R=>rst);
   ix20632 : oai21 port map ( Y=>nx20631, A0=>nx33152, A1=>nx42375, B0=>
      nx33154);
   booth_booth_integrtaion_0_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_25, QB=>nx33152, D=>nx20631, CLK=>clk, 
      R=>rst);
   ix33155 : nand03 port map ( Y=>nx33154, A0=>nx42381, A1=>nx2616, A2=>
      nx42377);
   ix2617 : xnor2 port map ( Y=>nx2616, A0=>nx33157, A1=>nx18207);
   ix33158 : aoi22 port map ( Y=>nx33157, A0=>
      booth_booth_integration_output_0_25, A1=>nx2420, B0=>nx2400, B1=>
      nx18205);
   ix2411 : nor02_2x port map ( Y=>nx2410, A0=>data_in(9), A1=>nx33145);
   ix33170 : xnor2 port map ( Y=>nx33169, A0=>nx2448, A1=>nx18209);
   ix2449 : oai22 port map ( Y=>nx2448, A0=>nx33157, A1=>nx33172, B0=>
      nx33181, B1=>nx42393);
   ix33175 : aoi32 port map ( Y=>nx33174, A0=>nx2430, A1=>nx41789, A2=>
      nx33179, B0=>data_in(10), B1=>nx41785);
   ix2431 : nand02 port map ( Y=>nx2430, A0=>nx33177, A1=>data_in(10));
   ix33180 : nand02 port map ( Y=>nx33179, A0=>nx32498, A1=>nx2410);
   booth_booth_integrtaion_0_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_26, QB=>nx33181, D=>nx20621, CLK=>clk, 
      R=>rst);
   ix20612 : oai21 port map ( Y=>nx20611, A0=>nx33186, A1=>nx42375, B0=>
      nx33188);
   booth_booth_integrtaion_0_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_27, QB=>nx33186, D=>nx20611, CLK=>clk, 
      R=>rst);
   ix33189 : nand03 port map ( Y=>nx33188, A0=>nx43131, A1=>nx2592, A2=>
      nx42377);
   ix2593 : xnor2 port map ( Y=>nx2592, A0=>nx33191, A1=>nx18210);
   ix33192 : aoi22 port map ( Y=>nx33191, A0=>
      booth_booth_integration_output_0_27, A1=>nx2468, B0=>nx2448, B1=>
      nx18209);
   ix2459 : nor02_2x port map ( Y=>nx2458, A0=>data_in(11), A1=>nx33179);
   ix33204 : xnor2 port map ( Y=>nx33203, A0=>nx2496, A1=>nx18211);
   ix2497 : oai22 port map ( Y=>nx2496, A0=>nx33191, A1=>nx33206, B0=>
      nx33215, B1=>nx42395);
   ix33209 : aoi32 port map ( Y=>nx33208, A0=>nx2478, A1=>nx41791, A2=>
      nx33213, B0=>data_in(12), B1=>nx41785);
   ix2479 : nand02 port map ( Y=>nx2478, A0=>nx33211, A1=>data_in(12));
   ix33214 : nand02 port map ( Y=>nx33213, A0=>nx32572, A1=>nx2458);
   booth_booth_integrtaion_0_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28, QB=>nx33215, D=>nx20601, CLK=>clk, R=>rst);
   ix20592 : oai21 port map ( Y=>nx20591, A0=>nx33220, A1=>nx42375, B0=>
      nx33222);
   booth_booth_integrtaion_0_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29, QB=>nx33220, D=>nx20591, CLK=>clk, R=>rst);
   ix33223 : nand03 port map ( Y=>nx33222, A0=>nx43131, A1=>nx2568, A2=>
      nx42375);
   ix2569 : xnor2 port map ( Y=>nx2568, A0=>nx33225, A1=>nx18212);
   ix33226 : aoi22 port map ( Y=>nx33225, A0=>booth_output_29, A1=>nx2516, 
      B0=>nx2496, B1=>nx18211);
   ix2507 : nor02_2x port map ( Y=>nx2506, A0=>data_in(13), A1=>nx33213);
   ix20582 : oai21 port map ( Y=>nx20581, A0=>nx33236, A1=>nx42375, B0=>
      nx33238);
   booth_booth_integrtaion_0_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx33236, D=>nx20581, CLK=>clk, R=>rst);
   ix33239 : nand03 port map ( Y=>nx33238, A0=>nx43131, A1=>nx2556, A2=>
      nx42375);
   ix2557 : xnor2 port map ( Y=>nx2556, A0=>nx2544, A1=>nx33251);
   ix2545 : oai22 port map ( Y=>nx2544, A0=>nx33225, A1=>nx33242, B0=>
      nx33236, B1=>nx42397);
   ix33245 : aoi32 port map ( Y=>nx33244, A0=>nx2526, A1=>nx41791, A2=>
      nx33249, B0=>data_in(14), B1=>nx41787);
   ix2527 : nand02 port map ( Y=>nx2526, A0=>nx33247, A1=>data_in(14));
   ix33250 : nand02 port map ( Y=>nx33249, A0=>nx32647, A1=>nx2506);
   ix2553 : oai22 port map ( Y=>nx2552, A0=>nx33023, A1=>nx33254, B0=>
      nx33256, B1=>nx33026);
   ix33255 : xnor2 port map ( Y=>nx33254, A0=>data_in(15), A1=>nx33249);
   ix33257 : inv01 port map ( Y=>nx33256, A=>data_in(15));
   ix33259 : aoi32 port map ( Y=>nx33258, A0=>nx2502, A1=>nx41791, A2=>
      nx33247, B0=>data_in(13), B1=>nx41787);
   ix2503 : nand02 port map ( Y=>nx2502, A0=>nx33213, A1=>data_in(13));
   ix33262 : aoi32 port map ( Y=>nx33261, A0=>nx2454, A1=>nx41791, A2=>
      nx33211, B0=>data_in(11), B1=>nx41787);
   ix2455 : nand02 port map ( Y=>nx2454, A0=>nx33179, A1=>data_in(11));
   ix33265 : aoi32 port map ( Y=>nx33264, A0=>nx2406, A1=>nx41791, A2=>
      nx33177, B0=>data_in(9), B1=>nx41787);
   ix2407 : nand02 port map ( Y=>nx2406, A0=>nx33145, A1=>data_in(9));
   ix33268 : aoi32 port map ( Y=>nx33267, A0=>nx2358, A1=>nx41791, A2=>
      nx33143, B0=>data_in(7), B1=>nx41787);
   ix2359 : nand02 port map ( Y=>nx2358, A0=>nx33111, A1=>data_in(7));
   ix33271 : aoi32 port map ( Y=>nx33270, A0=>nx2310, A1=>nx41793, A2=>
      nx33109, B0=>data_in(5), B1=>nx41787);
   ix2311 : nand02 port map ( Y=>nx2310, A0=>nx33077, A1=>data_in(5));
   ix33274 : aoi32 port map ( Y=>nx33273, A0=>nx2212, A1=>nx41793, A2=>
      nx33276, B0=>data_in(1), B1=>nx41787);
   ix2213 : nand02 port map ( Y=>nx2212, A0=>data_in(1), A1=>data_in(0));
   booth_booth_integrtaion_0_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_16, QB=>nx33001, D=>nx20721, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_15, QB=>nx33280, D=>nx20741, CLK=>clk, 
      R=>rst);
   reg_neuron_14 : dff port map ( Q=>neuron_14, QB=>OPEN, D=>nx20751, CLK=>
      clk);
   reg_neuron_13 : dff port map ( Q=>neuron_13, QB=>OPEN, D=>nx20771, CLK=>
      clk);
   reg_neuron_12 : dff port map ( Q=>neuron_12, QB=>OPEN, D=>nx20791, CLK=>
      clk);
   ix2819 : aoi21 port map ( Y=>nx2818, A0=>label_1_output_0, A1=>
      booth_booth_integration_output_0_12, B0=>nx43519);
   reg_sel_dst_0 : dffr port map ( Q=>sel_dst_0, QB=>OPEN, D=>nx20111, CLK=>
      clk, R=>rst);
   ix20112 : mux21_ni port map ( Y=>nx20111, A0=>sel_dst_0, A1=>nx43349, S0
      =>nx1860);
   ix1861 : aoi321 port map ( Y=>nx1860, A0=>nx33302, A1=>nx33304, A2=>
      nx42865, B0=>nx122, B1=>nx41379, C0=>nx104);
   ix33303 : nand02 port map ( Y=>nx33302, A0=>nx33299, A1=>nx31961);
   ix33305 : oai221 port map ( Y=>nx33304, A0=>nx41397, A1=>nx42891, B0=>
      nx43103, B1=>nx31961, C0=>nx36);
   labelsregfile_label1_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_1_output_1, QB=>nx33325, D=>nx30131, CLK=>clk, R=>rst);
   lat_label_1_input_1 : latch port map ( Q=>label_1_input_1, D=>nx17648, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_1 : dffr port map ( Q=>
      label_1_input_state_machine_1, QB=>OPEN, D=>nx30121, CLK=>clk, R=>rst
   );
   ix17645 : xor2 port map ( Y=>nx17644, A0=>nx32810, A1=>nx33315);
   ix33327 : xnor2 port map ( Y=>nx33326, A0=>
      booth_booth_integration_output_0_14, A1=>label_1_output_2);
   labelsregfile_label1_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_1_output_3, QB=>nx33340, D=>nx30171, CLK=>clk, R=>rst);
   lat_label_1_input_3 : latch port map ( Q=>label_1_input_3, D=>nx17712, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_3 : dffr port map ( Q=>
      label_1_input_state_machine_3, QB=>OPEN, D=>nx30161, CLK=>clk, R=>rst
   );
   ix17709 : xor2 port map ( Y=>nx17708, A0=>nx32799, A1=>nx33330);
   labelsregfile_label1_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_1_output_5, QB=>nx33355, D=>nx30211, CLK=>clk, R=>rst);
   lat_label_1_input_5 : latch port map ( Q=>label_1_input_5, D=>nx17776, 
      CLK=>nx41661);
   reg_label_1_input_state_machine_5 : dffr port map ( Q=>
      label_1_input_state_machine_5, QB=>OPEN, D=>nx30201, CLK=>clk, R=>rst
   );
   ix17773 : xor2 port map ( Y=>nx17772, A0=>nx32788, A1=>nx33345);
   labelsregfile_label1_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_1_output_7, QB=>nx33370, D=>nx30251, CLK=>clk, R=>rst);
   lat_label_1_input_7 : latch port map ( Q=>label_1_input_7, D=>nx17840, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_7 : dffr port map ( Q=>
      label_1_input_state_machine_7, QB=>OPEN, D=>nx30241, CLK=>clk, R=>rst
   );
   ix17837 : xor2 port map ( Y=>nx17836, A0=>nx32777, A1=>nx33360);
   labelsregfile_label1_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_1_output_9, QB=>nx33385, D=>nx30291, CLK=>clk, R=>rst);
   lat_label_1_input_9 : latch port map ( Q=>label_1_input_9, D=>nx17904, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_9 : dffr port map ( Q=>
      label_1_input_state_machine_9, QB=>OPEN, D=>nx30281, CLK=>clk, R=>rst
   );
   ix17901 : xor2 port map ( Y=>nx17900, A0=>nx32766, A1=>nx33375);
   labelsregfile_label1_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_1_output_11, QB=>nx33400, D=>nx30331, CLK=>clk, R=>rst);
   lat_label_1_input_11 : latch port map ( Q=>label_1_input_11, D=>nx17968, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_11 : dffr port map ( Q=>
      label_1_input_state_machine_11, QB=>OPEN, D=>nx30321, CLK=>clk, R=>rst
   );
   ix17965 : xor2 port map ( Y=>nx17964, A0=>nx32755, A1=>nx33390);
   labelsregfile_label1_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_1_output_13, QB=>nx33415, D=>nx30371, CLK=>clk, R=>rst);
   lat_label_1_input_13 : latch port map ( Q=>label_1_input_13, D=>nx18032, 
      CLK=>nx41663);
   reg_label_1_input_state_machine_13 : dffr port map ( Q=>
      label_1_input_state_machine_13, QB=>OPEN, D=>nx30361, CLK=>clk, R=>rst
   );
   ix18029 : xor2 port map ( Y=>nx18028, A0=>nx32744, A1=>nx33405);
   labelsregfile_label1_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_1_output_15, QB=>nx33421, D=>nx31581, CLK=>clk, R=>rst);
   max_calc_reg_ans1_15 : dff port map ( Q=>max_calc_ans1_15, QB=>OPEN, D=>
      nx31591, CLK=>clk);
   max_calc_reg_state_2 : dffr port map ( Q=>max_calc_state_2, QB=>OPEN, D=>
      nx20081, CLK=>clk, R=>rst);
   ix31822 : oai21 port map ( Y=>nx31821, A0=>nx42925, A1=>nx1714, B0=>
      nx33432);
   max_calc_reg_state_3 : dffr port map ( Q=>OPEN, QB=>nx33429, D=>nx31821, 
      CLK=>clk, R=>rst);
   ix33433 : oai21 port map ( Y=>nx33432, A0=>nx20920, A1=>nx18191, B0=>
      max_calc_start);
   ix20921 : oai21 port map ( Y=>nx20920, A0=>nx18189, A1=>nx18187, B0=>
      nx41577);
   max_calc_reg_state_0 : dffr port map ( Q=>max_calc_state_0, QB=>nx33436, 
      D=>nx20091, CLK=>clk, R=>rst);
   ix20102 : ao32 port map ( Y=>nx20101, A0=>nx18183, A1=>nx42925, A2=>
      max_calc_start, B0=>nx41535, B1=>nx33444);
   ix1791 : oai21 port map ( Y=>nx18183, A0=>max_calc_state_0, A1=>nx43137, 
      B0=>nx1782);
   max_calc_reg_state_1 : dffr port map ( Q=>max_calc_state_1, QB=>OPEN, D=>
      nx20101, CLK=>clk, R=>rst);
   ix20911 : nor04 port map ( Y=>nx18191, A0=>nx20772, A1=>nx33450, A2=>
      nx40947, A3=>nx40985);
   ix33451 : nor04 port map ( Y=>nx33450, A0=>nx20830, A1=>nx20816, A2=>
      nx20800, A3=>nx20786);
   ix20831 : nand04 port map ( Y=>nx20830, A0=>nx33453, A1=>nx34097, A2=>
      nx40874, A3=>nx40879);
   lat_label_10_input_15 : latch port map ( Q=>label_10_input_15, D=>nx5916, 
      CLK=>nx41669);
   reg_label_10_input_state_machine_15 : dffr port map ( Q=>
      label_10_input_state_machine_15, QB=>OPEN, D=>nx22811, CLK=>clk, R=>
      rst);
   ix5913 : xnor2 port map ( Y=>nx5912, A0=>nx33463, A1=>nx5910);
   ix33464 : aoi22 port map ( Y=>nx33463, A0=>label_10_output_14, A1=>
      booth_booth_integration_output_9_26, B0=>nx5054, B1=>nx5056);
   labelsregfile_label10_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_10_output_14, QB=>OPEN, D=>nx22231, CLK=>clk, R=>rst);
   lat_label_10_input_14 : latch port map ( Q=>label_10_input_14, D=>nx5062, 
      CLK=>nx41669);
   reg_label_10_input_state_machine_14 : dffr port map ( Q=>
      label_10_input_state_machine_14, QB=>OPEN, D=>nx21411, CLK=>clk, R=>
      rst);
   ix5059 : xnor2 port map ( Y=>nx5058, A0=>nx5054, A1=>nx34090);
   ix5055 : oai22 port map ( Y=>nx5054, A0=>nx33474, A1=>nx34079, B0=>
      nx34089, B1=>nx33848);
   ix33475 : aoi22 port map ( Y=>nx33474, A0=>label_10_output_12, A1=>
      booth_booth_integration_output_9_24, B0=>nx4990, B1=>nx18271);
   labelsregfile_label10_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_10_output_12, QB=>OPEN, D=>nx22201, CLK=>clk, R=>rst);
   lat_label_10_input_12 : latch port map ( Q=>label_10_input_12, D=>nx5004, 
      CLK=>nx41669);
   reg_label_10_input_state_machine_12 : dffr port map ( Q=>
      label_10_input_state_machine_12, QB=>OPEN, D=>nx22191, CLK=>clk, R=>
      rst);
   ix5001 : xnor2 port map ( Y=>nx5000, A0=>nx4990, A1=>nx34075);
   ix4991 : oai22 port map ( Y=>nx4990, A0=>nx33485, A1=>nx34064, B0=>
      nx34074, B1=>nx33812);
   ix33486 : aoi22 port map ( Y=>nx33485, A0=>label_10_output_10, A1=>
      booth_booth_integration_output_9_22, B0=>nx4926, B1=>nx18268);
   labelsregfile_label10_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_10_output_10, QB=>OPEN, D=>nx22161, CLK=>clk, R=>rst);
   lat_label_10_input_10 : latch port map ( Q=>label_10_input_10, D=>nx4940, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_10 : dffr port map ( Q=>
      label_10_input_state_machine_10, QB=>OPEN, D=>nx22151, CLK=>clk, R=>
      rst);
   ix4937 : xnor2 port map ( Y=>nx4936, A0=>nx4926, A1=>nx34060);
   ix4927 : oai22 port map ( Y=>nx4926, A0=>nx33496, A1=>nx34049, B0=>
      nx34059, B1=>nx33776);
   ix33497 : aoi22 port map ( Y=>nx33496, A0=>label_10_output_8, A1=>
      booth_booth_integration_output_9_20, B0=>nx4862, B1=>nx18266);
   labelsregfile_label10_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_10_output_8, QB=>OPEN, D=>nx22121, CLK=>clk, R=>rst);
   lat_label_10_input_8 : latch port map ( Q=>label_10_input_8, D=>nx4876, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_8 : dffr port map ( Q=>
      label_10_input_state_machine_8, QB=>OPEN, D=>nx22111, CLK=>clk, R=>rst
   );
   ix4873 : xnor2 port map ( Y=>nx4872, A0=>nx4862, A1=>nx34045);
   ix4863 : oai22 port map ( Y=>nx4862, A0=>nx33507, A1=>nx34034, B0=>
      nx34044, B1=>nx33738);
   ix33508 : aoi22 port map ( Y=>nx33507, A0=>label_10_output_6, A1=>
      booth_booth_integration_output_9_18, B0=>nx4798, B1=>nx18264);
   labelsregfile_label10_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_10_output_6, QB=>OPEN, D=>nx22081, CLK=>clk, R=>rst);
   lat_label_10_input_6 : latch port map ( Q=>label_10_input_6, D=>nx4812, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_6 : dffr port map ( Q=>
      label_10_input_state_machine_6, QB=>OPEN, D=>nx22071, CLK=>clk, R=>rst
   );
   ix4809 : xnor2 port map ( Y=>nx4808, A0=>nx4798, A1=>nx34030);
   ix4799 : oai22 port map ( Y=>nx4798, A0=>nx33518, A1=>nx34019, B0=>
      nx34029, B1=>nx33699);
   ix33519 : aoi22 port map ( Y=>nx33518, A0=>label_10_output_4, A1=>
      booth_booth_integration_output_9_16, B0=>nx4734, B1=>nx18261);
   labelsregfile_label10_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_10_output_4, QB=>OPEN, D=>nx22041, CLK=>clk, R=>rst);
   lat_label_10_input_4 : latch port map ( Q=>label_10_input_4, D=>nx4748, 
      CLK=>nx41665);
   reg_label_10_input_state_machine_4 : dffr port map ( Q=>
      label_10_input_state_machine_4, QB=>OPEN, D=>nx22031, CLK=>clk, R=>rst
   );
   ix4745 : xnor2 port map ( Y=>nx4744, A0=>nx4734, A1=>nx34015);
   ix4735 : oai22 port map ( Y=>nx4734, A0=>nx33529, A1=>nx34004, B0=>
      nx34014, B1=>nx33982);
   ix33530 : aoi22 port map ( Y=>nx33529, A0=>label_10_output_2, A1=>
      booth_booth_integration_output_9_14, B0=>nx4670, B1=>nx18259);
   labelsregfile_label10_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_10_output_2, QB=>OPEN, D=>nx22001, CLK=>clk, R=>rst);
   lat_label_10_input_2 : latch port map ( Q=>label_10_input_2, D=>nx4684, 
      CLK=>nx41665);
   reg_label_10_input_state_machine_2 : dffr port map ( Q=>
      label_10_input_state_machine_2, QB=>OPEN, D=>nx21991, CLK=>clk, R=>rst
   );
   ix4681 : xnor2 port map ( Y=>nx4680, A0=>nx4670, A1=>nx34000);
   ix4671 : oai22 port map ( Y=>nx4670, A0=>nx33540, A1=>nx33989, B0=>
      nx33999, B1=>nx33985);
   ix33541 : nand02 port map ( Y=>nx33540, A0=>label_10_output_0, A1=>
      booth_booth_integration_output_9_12);
   labelsregfile_label10_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_10_output_0, QB=>OPEN, D=>nx21961, CLK=>clk, R=>rst);
   lat_label_10_input_0 : latch port map ( Q=>label_10_input_0, D=>nx4626, 
      CLK=>nx41665);
   ix4627 : oai21 port map ( Y=>nx4626, A0=>nx33546, A1=>nx41425, B0=>
      nx33550);
   reg_label_10_input_state_machine_0 : dffr port map ( Q=>
      label_10_input_state_machine_0, QB=>nx33546, D=>nx21951, CLK=>clk, R=>
      rst);
   ix33551 : oai21 port map ( Y=>nx33550, A0=>
      booth_booth_integration_output_9_12, A1=>label_10_output_0, B0=>nx4614
   );
   booth_booth_integrtaion_9_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_12, QB=>OPEN, D=>nx21941, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_13, QB=>nx33985, D=>nx21931, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_14, QB=>OPEN, D=>nx21921, CLK=>clk, R
      =>rst);
   ix33564 : aoi22 port map ( Y=>nx33563, A0=>nx41795, A1=>nx41879, B0=>
      nx4556, B1=>nx4562);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_reg_output_0, QB=>OPEN, 
      D=>nx21441, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_0, QB=>OPEN, D=>nx21427, CLK
      =>clk, S=>nx41481);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_reg_output_9, QB=>OPEN, 
      D=>nx21621, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_9, QB=>OPEN, D=>nx21611, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12940, QB=>OPEN, D=>nx21601, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_8, QB=>OPEN, D=>nx21591, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12941, QB=>OPEN, D=>nx21581, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_7, QB=>OPEN, D=>nx21571, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12942, QB=>OPEN, D=>nx21561, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_6, QB=>OPEN, D=>nx21551, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12943, QB=>OPEN, D=>nx21541, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_5, QB=>OPEN, D=>nx21531, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12944, QB=>OPEN, D=>nx21521, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_4, QB=>OPEN, D=>nx21511, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12945, QB=>OPEN, D=>nx21501, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_3, QB=>OPEN, D=>nx21491, CLK
      =>clk, R=>nx41479);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12946, QB=>OPEN, D=>nx21481, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_2, QB=>OPEN, D=>nx21471, CLK
      =>clk, R=>nx41477);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12947, QB=>OPEN, D=>nx21461, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_1, QB=>OPEN, D=>nx21451, CLK
      =>clk, R=>nx41477);
   ix21422 : nand02 port map ( Y=>nx21421, A0=>nx42929, A1=>nx41865);
   booth_booth_integrtaion_9_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx33610, D=>nx21421, CLK=>clk, S=>nx41477);
   ix4557 : nand02 port map ( Y=>nx4556, A0=>nx33631, A1=>nx33689);
   ix33632 : oai21 port map ( Y=>nx33631, A0=>nx41891, A1=>nx41887, B0=>
      data_in(144));
   ix21752 : oai21 port map ( Y=>nx21751, A0=>nx33636, A1=>nx42459, B0=>
      nx33638);
   booth_booth_integrtaion_9_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx33636, D=>nx21751, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12282, QB=>nx33687, D=>nx21741, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12281, QB=>OPEN, D=>nx21731, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12280, QB=>OPEN, D=>nx21721, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12279, QB=>OPEN, D=>nx21711, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12278, QB=>OPEN, D=>nx21701, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12277, QB=>OPEN, D=>nx21691, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12276, QB=>OPEN, D=>nx21681, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12275, QB=>OPEN, D=>nx21671, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12274, QB=>OPEN, D=>nx21661, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12273, QB=>OPEN, D=>nx21651, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12272, QB=>OPEN, D=>nx21641, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12271, QB=>OPEN, D=>nx21631, CLK=>clk, R=>rst);
   ix33694 : xnor2 port map ( Y=>nx33693, A0=>nx4026, A1=>nx18239);
   ix21892 : oai21 port map ( Y=>nx21891, A0=>nx33699, A1=>nx42459, B0=>
      nx33701);
   booth_booth_integrtaion_9_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_17, QB=>nx33699, D=>nx21891, CLK=>clk, 
      R=>rst);
   ix33702 : nand03 port map ( Y=>nx33701, A0=>nx42467, A1=>nx4534, A2=>
      nx42463);
   ix4535 : xnor2 port map ( Y=>nx4534, A0=>nx33704, A1=>nx18241);
   ix33705 : aoi22 port map ( Y=>nx33704, A0=>
      booth_booth_integration_output_9_17, A1=>nx4050, B0=>nx4026, B1=>
      nx18239);
   ix4041 : nor02_2x port map ( Y=>nx4040, A0=>data_in(144), A1=>
      data_in(145));
   ix21882 : oai21 port map ( Y=>nx21881, A0=>nx33719, A1=>nx42459, B0=>
      nx33721);
   booth_booth_integrtaion_9_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_18, QB=>nx33719, D=>nx21881, CLK=>clk, 
      R=>rst);
   ix33722 : nand03 port map ( Y=>nx33721, A0=>nx42467, A1=>nx4522, A2=>
      nx42463);
   ix4523 : xnor2 port map ( Y=>nx4522, A0=>nx4078, A1=>nx33734);
   ix4079 : oai22 port map ( Y=>nx4078, A0=>nx33704, A1=>nx33725, B0=>
      nx33719, B1=>nx42471);
   ix33728 : aoi32 port map ( Y=>nx33727, A0=>nx4060, A1=>nx41891, A2=>
      nx33730, B0=>data_in(146), B1=>nx41887);
   ix4061 : oai21 port map ( Y=>nx4060, A0=>data_in(144), A1=>data_in(145), 
      B0=>data_in(146));
   ix21872 : oai21 port map ( Y=>nx21871, A0=>nx33738, A1=>nx42459, B0=>
      nx33740);
   booth_booth_integrtaion_9_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_19, QB=>nx33738, D=>nx21871, CLK=>clk, 
      R=>rst);
   ix33741 : nand03 port map ( Y=>nx33740, A0=>nx42467, A1=>nx4510, A2=>
      nx42463);
   ix4511 : xnor2 port map ( Y=>nx4510, A0=>nx33743, A1=>nx18243);
   ix33744 : aoi22 port map ( Y=>nx33743, A0=>
      booth_booth_integration_output_9_19, A1=>nx4098, B0=>nx4078, B1=>
      nx18242);
   ix4099 : oai32 port map ( Y=>nx4098, A0=>nx33746, A1=>nx33709, A2=>nx4088, 
      B0=>nx33749, B1=>nx33714);
   ix4065 : nor03_2x port map ( Y=>nx4064, A0=>data_in(146), A1=>
      data_in(144), A2=>data_in(145));
   ix33750 : inv01 port map ( Y=>nx33749, A=>data_in(147));
   ix4089 : nor04 port map ( Y=>nx4088, A0=>data_in(147), A1=>data_in(146), 
      A2=>data_in(144), A3=>data_in(145));
   ix33758 : xnor2 port map ( Y=>nx33757, A0=>nx4126, A1=>nx18244);
   ix4127 : oai22 port map ( Y=>nx4126, A0=>nx33743, A1=>nx33760, B0=>
      nx33771, B1=>nx42473);
   ix33763 : aoi32 port map ( Y=>nx33762, A0=>nx4108, A1=>nx41891, A2=>
      nx33767, B0=>data_in(148), B1=>nx41887);
   ix4109 : nand02 port map ( Y=>nx4108, A0=>nx33765, A1=>data_in(148));
   ix33768 : nand02 port map ( Y=>nx33767, A0=>nx33769, A1=>nx4088);
   ix33770 : inv01 port map ( Y=>nx33769, A=>data_in(148));
   booth_booth_integrtaion_9_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_20, QB=>nx33771, D=>nx21861, CLK=>clk, 
      R=>rst);
   ix21852 : oai21 port map ( Y=>nx21851, A0=>nx33776, A1=>nx42459, B0=>
      nx33778);
   booth_booth_integrtaion_9_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_21, QB=>nx33776, D=>nx21851, CLK=>clk, 
      R=>rst);
   ix33779 : nand03 port map ( Y=>nx33778, A0=>nx42467, A1=>nx4486, A2=>
      nx42463);
   ix4487 : xnor2 port map ( Y=>nx4486, A0=>nx33781, A1=>nx18245);
   ix33782 : aoi22 port map ( Y=>nx33781, A0=>
      booth_booth_integration_output_9_21, A1=>nx4146, B0=>nx4126, B1=>
      nx18244);
   ix4137 : nor02_2x port map ( Y=>nx4136, A0=>data_in(149), A1=>nx33767);
   ix33794 : xnor2 port map ( Y=>nx33793, A0=>nx4174, A1=>nx18246);
   ix4175 : oai22 port map ( Y=>nx4174, A0=>nx33781, A1=>nx33796, B0=>
      nx33807, B1=>nx42475);
   ix33799 : aoi32 port map ( Y=>nx33798, A0=>nx4156, A1=>nx41891, A2=>
      nx33803, B0=>data_in(150), B1=>nx41887);
   ix4157 : nand02 port map ( Y=>nx4156, A0=>nx33801, A1=>data_in(150));
   ix33804 : nand02 port map ( Y=>nx33803, A0=>nx33805, A1=>nx4136);
   ix33806 : inv01 port map ( Y=>nx33805, A=>data_in(150));
   booth_booth_integrtaion_9_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_22, QB=>nx33807, D=>nx21841, CLK=>clk, 
      R=>rst);
   ix21832 : oai21 port map ( Y=>nx21831, A0=>nx33812, A1=>nx42461, B0=>
      nx33814);
   booth_booth_integrtaion_9_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_23, QB=>nx33812, D=>nx21831, CLK=>clk, 
      R=>rst);
   ix33815 : nand03 port map ( Y=>nx33814, A0=>nx42467, A1=>nx4462, A2=>
      nx42463);
   ix4463 : xnor2 port map ( Y=>nx4462, A0=>nx33817, A1=>nx18247);
   ix33818 : aoi22 port map ( Y=>nx33817, A0=>
      booth_booth_integration_output_9_23, A1=>nx4194, B0=>nx4174, B1=>
      nx18246);
   ix4185 : nor02_2x port map ( Y=>nx4184, A0=>data_in(151), A1=>nx33803);
   ix33830 : xnor2 port map ( Y=>nx33829, A0=>nx4222, A1=>nx18249);
   ix4223 : oai22 port map ( Y=>nx4222, A0=>nx33817, A1=>nx33832, B0=>
      nx33843, B1=>nx42477);
   ix33835 : aoi32 port map ( Y=>nx33834, A0=>nx4204, A1=>nx41891, A2=>
      nx33839, B0=>data_in(152), B1=>nx41887);
   ix4205 : nand02 port map ( Y=>nx4204, A0=>nx33837, A1=>data_in(152));
   ix33840 : nand02 port map ( Y=>nx33839, A0=>nx33841, A1=>nx4184);
   ix33842 : inv01 port map ( Y=>nx33841, A=>data_in(152));
   booth_booth_integrtaion_9_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_24, QB=>nx33843, D=>nx21821, CLK=>clk, 
      R=>rst);
   ix21812 : oai21 port map ( Y=>nx21811, A0=>nx33848, A1=>nx42461, B0=>
      nx33850);
   booth_booth_integrtaion_9_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_25, QB=>nx33848, D=>nx21811, CLK=>clk, 
      R=>rst);
   ix33851 : nand03 port map ( Y=>nx33850, A0=>nx42467, A1=>nx4438, A2=>
      nx42463);
   ix4439 : xnor2 port map ( Y=>nx4438, A0=>nx33853, A1=>nx18251);
   ix33854 : aoi22 port map ( Y=>nx33853, A0=>
      booth_booth_integration_output_9_25, A1=>nx4242, B0=>nx4222, B1=>
      nx18249);
   ix4233 : nor02_2x port map ( Y=>nx4232, A0=>data_in(153), A1=>nx33839);
   ix33866 : xnor2 port map ( Y=>nx33865, A0=>nx4270, A1=>nx18253);
   ix4271 : oai22 port map ( Y=>nx4270, A0=>nx33853, A1=>nx33868, B0=>
      nx33879, B1=>nx42479);
   ix33871 : aoi32 port map ( Y=>nx33870, A0=>nx4252, A1=>nx41891, A2=>
      nx33875, B0=>data_in(154), B1=>nx41887);
   ix4253 : nand02 port map ( Y=>nx4252, A0=>nx33873, A1=>data_in(154));
   ix33876 : nand02 port map ( Y=>nx33875, A0=>nx33877, A1=>nx4232);
   ix33878 : inv01 port map ( Y=>nx33877, A=>data_in(154));
   booth_booth_integrtaion_9_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_26, QB=>nx33879, D=>nx21801, CLK=>clk, 
      R=>rst);
   ix21792 : oai21 port map ( Y=>nx21791, A0=>nx33884, A1=>nx42461, B0=>
      nx33886);
   booth_booth_integrtaion_9_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_27, QB=>nx33884, D=>nx21791, CLK=>clk, 
      R=>rst);
   ix33887 : nand03 port map ( Y=>nx33886, A0=>nx43171, A1=>nx4414, A2=>
      nx42463);
   ix4415 : xnor2 port map ( Y=>nx4414, A0=>nx33889, A1=>nx18254);
   ix33890 : aoi22 port map ( Y=>nx33889, A0=>
      booth_booth_integration_output_9_27, A1=>nx4290, B0=>nx4270, B1=>
      nx18253);
   ix4281 : nor02_2x port map ( Y=>nx4280, A0=>data_in(155), A1=>nx33875);
   ix33902 : xnor2 port map ( Y=>nx33901, A0=>nx4318, A1=>nx18255);
   ix4319 : oai22 port map ( Y=>nx4318, A0=>nx33889, A1=>nx33904, B0=>
      nx33915, B1=>nx42481);
   ix33907 : aoi32 port map ( Y=>nx33906, A0=>nx4300, A1=>nx41893, A2=>
      nx33911, B0=>data_in(156), B1=>nx41887);
   ix4301 : nand02 port map ( Y=>nx4300, A0=>nx33909, A1=>data_in(156));
   ix33912 : nand02 port map ( Y=>nx33911, A0=>nx33913, A1=>nx4280);
   ix33914 : inv01 port map ( Y=>nx33913, A=>data_in(156));
   booth_booth_integrtaion_9_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12270, QB=>nx33915, D=>nx21781, CLK=>clk, R=>rst);
   ix21772 : oai21 port map ( Y=>nx21771, A0=>nx33920, A1=>nx42461, B0=>
      nx33922);
   booth_booth_integrtaion_9_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12269, QB=>nx33920, D=>nx21771, CLK=>clk, R=>rst);
   ix33923 : nand03 port map ( Y=>nx33922, A0=>nx43171, A1=>nx4390, A2=>
      nx42461);
   ix4391 : xnor2 port map ( Y=>nx4390, A0=>nx33925, A1=>nx18256);
   ix33926 : aoi22 port map ( Y=>nx33925, A0=>booth_output_29_dup_12269, A1
      =>nx4338, B0=>nx4318, B1=>nx18255);
   ix4329 : nor02_2x port map ( Y=>nx4328, A0=>data_in(157), A1=>nx33911);
   ix21762 : oai21 port map ( Y=>nx21761, A0=>nx33936, A1=>nx42461, B0=>
      nx33938);
   booth_booth_integrtaion_9_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx33936, D=>nx21761, CLK=>clk, R=>rst);
   ix33939 : nand03 port map ( Y=>nx33938, A0=>nx43171, A1=>nx4378, A2=>
      nx42461);
   ix4379 : xnor2 port map ( Y=>nx4378, A0=>nx4366, A1=>nx33953);
   ix4367 : oai22 port map ( Y=>nx4366, A0=>nx33925, A1=>nx33942, B0=>
      nx33936, B1=>nx42483);
   ix33945 : aoi32 port map ( Y=>nx33944, A0=>nx4348, A1=>nx41893, A2=>
      nx33949, B0=>data_in(158), B1=>nx41889);
   ix4349 : nand02 port map ( Y=>nx4348, A0=>nx33947, A1=>data_in(158));
   ix33950 : nand02 port map ( Y=>nx33949, A0=>nx33951, A1=>nx4328);
   ix33952 : inv01 port map ( Y=>nx33951, A=>data_in(158));
   ix4375 : oai22 port map ( Y=>nx4374, A0=>nx33709, A1=>nx33956, B0=>
      nx33958, B1=>nx33714);
   ix33957 : xnor2 port map ( Y=>nx33956, A0=>data_in(159), A1=>nx33949);
   ix33959 : inv01 port map ( Y=>nx33958, A=>data_in(159));
   ix33961 : aoi32 port map ( Y=>nx33960, A0=>nx4324, A1=>nx41893, A2=>
      nx33947, B0=>data_in(157), B1=>nx41889);
   ix4325 : nand02 port map ( Y=>nx4324, A0=>nx33911, A1=>data_in(157));
   ix33964 : aoi32 port map ( Y=>nx33963, A0=>nx4276, A1=>nx41893, A2=>
      nx33909, B0=>data_in(155), B1=>nx41889);
   ix4277 : nand02 port map ( Y=>nx4276, A0=>nx33875, A1=>data_in(155));
   ix33967 : aoi32 port map ( Y=>nx33966, A0=>nx4228, A1=>nx41893, A2=>
      nx33873, B0=>data_in(153), B1=>nx41889);
   ix4229 : nand02 port map ( Y=>nx4228, A0=>nx33839, A1=>data_in(153));
   ix33970 : aoi32 port map ( Y=>nx33969, A0=>nx4180, A1=>nx41893, A2=>
      nx33837, B0=>data_in(151), B1=>nx41889);
   ix4181 : nand02 port map ( Y=>nx4180, A0=>nx33803, A1=>data_in(151));
   ix33973 : aoi32 port map ( Y=>nx33972, A0=>nx4132, A1=>nx41895, A2=>
      nx33801, B0=>data_in(149), B1=>nx41889);
   ix4133 : nand02 port map ( Y=>nx4132, A0=>nx33767, A1=>data_in(149));
   ix33976 : aoi32 port map ( Y=>nx33975, A0=>nx4034, A1=>nx41895, A2=>
      nx33978, B0=>data_in(145), B1=>nx41889);
   ix4035 : nand02 port map ( Y=>nx4034, A0=>data_in(145), A1=>data_in(144)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_16, QB=>nx33689, D=>nx21901, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_15, QB=>nx33982, D=>nx21911, CLK=>clk, 
      R=>rst);
   ix4615 : aoi21 port map ( Y=>nx4614, A0=>label_10_output_0, A1=>
      booth_booth_integration_output_9_12, B0=>nx43519);
   labelsregfile_label10_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_10_output_1, QB=>nx33999, D=>nx21981, CLK=>clk, R=>rst);
   lat_label_10_input_1 : latch port map ( Q=>label_10_input_1, D=>nx4652, 
      CLK=>nx41665);
   reg_label_10_input_state_machine_1 : dffr port map ( Q=>
      label_10_input_state_machine_1, QB=>OPEN, D=>nx21971, CLK=>clk, R=>rst
   );
   ix4649 : xor2 port map ( Y=>nx4648, A0=>nx33540, A1=>nx33989);
   ix34001 : xnor2 port map ( Y=>nx34000, A0=>
      booth_booth_integration_output_9_14, A1=>label_10_output_2);
   labelsregfile_label10_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_10_output_3, QB=>nx34014, D=>nx22021, CLK=>clk, R=>rst);
   lat_label_10_input_3 : latch port map ( Q=>label_10_input_3, D=>nx4716, 
      CLK=>nx41665);
   reg_label_10_input_state_machine_3 : dffr port map ( Q=>
      label_10_input_state_machine_3, QB=>OPEN, D=>nx22011, CLK=>clk, R=>rst
   );
   ix4713 : xor2 port map ( Y=>nx4712, A0=>nx33529, A1=>nx34004);
   labelsregfile_label10_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_10_output_5, QB=>nx34029, D=>nx22061, CLK=>clk, R=>rst);
   lat_label_10_input_5 : latch port map ( Q=>label_10_input_5, D=>nx4780, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_5 : dffr port map ( Q=>
      label_10_input_state_machine_5, QB=>OPEN, D=>nx22051, CLK=>clk, R=>rst
   );
   ix4777 : xor2 port map ( Y=>nx4776, A0=>nx33518, A1=>nx34019);
   labelsregfile_label10_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_10_output_7, QB=>nx34044, D=>nx22101, CLK=>clk, R=>rst);
   lat_label_10_input_7 : latch port map ( Q=>label_10_input_7, D=>nx4844, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_7 : dffr port map ( Q=>
      label_10_input_state_machine_7, QB=>OPEN, D=>nx22091, CLK=>clk, R=>rst
   );
   ix4841 : xor2 port map ( Y=>nx4840, A0=>nx33507, A1=>nx34034);
   labelsregfile_label10_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_10_output_9, QB=>nx34059, D=>nx22141, CLK=>clk, R=>rst);
   lat_label_10_input_9 : latch port map ( Q=>label_10_input_9, D=>nx4908, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_9 : dffr port map ( Q=>
      label_10_input_state_machine_9, QB=>OPEN, D=>nx22131, CLK=>clk, R=>rst
   );
   ix4905 : xor2 port map ( Y=>nx4904, A0=>nx33496, A1=>nx34049);
   labelsregfile_label10_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_10_output_11, QB=>nx34074, D=>nx22181, CLK=>clk, R=>rst);
   lat_label_10_input_11 : latch port map ( Q=>label_10_input_11, D=>nx4972, 
      CLK=>nx41667);
   reg_label_10_input_state_machine_11 : dffr port map ( Q=>
      label_10_input_state_machine_11, QB=>OPEN, D=>nx22171, CLK=>clk, R=>
      rst);
   ix4969 : xor2 port map ( Y=>nx4968, A0=>nx33485, A1=>nx34064);
   labelsregfile_label10_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_10_output_13, QB=>nx34089, D=>nx22221, CLK=>clk, R=>rst);
   lat_label_10_input_13 : latch port map ( Q=>label_10_input_13, D=>nx5036, 
      CLK=>nx41669);
   reg_label_10_input_state_machine_13 : dffr port map ( Q=>
      label_10_input_state_machine_13, QB=>OPEN, D=>nx22211, CLK=>clk, R=>
      rst);
   ix5033 : xor2 port map ( Y=>nx5032, A0=>nx33474, A1=>nx34079);
   labelsregfile_label10_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_10_output_15, QB=>nx34095, D=>nx22821, CLK=>clk, R=>rst);
   ix34098 : xnor2 port map ( Y=>nx34097, A0=>nx42213, A1=>
      label_10_output_14);
   max_calc_reg_answer_14 : dffr port map ( Q=>max_calc_answer_14, QB=>OPEN, 
      D=>nx31801, CLK=>clk, R=>rst);
   max_calc_reg_comparator_first_inp1_14 : dff port map ( Q=>
      max_calc_comparator_first_inp1_14, QB=>OPEN, D=>nx30421, CLK=>clk);
   max_calc_reg_ans1_14 : dff port map ( Q=>max_calc_ans1_14, QB=>OPEN, D=>
      nx30391, CLK=>clk);
   max_calc_reg_ans6_14 : dff port map ( Q=>max_calc_ans6_14, QB=>OPEN, D=>
      nx30401, CLK=>clk);
   max_calc_reg_ans5_14 : dff port map ( Q=>max_calc_ans5_14, QB=>OPEN, D=>
      nx30411, CLK=>clk);
   ix22532 : oai21 port map ( Y=>nx22531, A0=>nx34125, A1=>nx41587, B0=>
      nx34128);
   max_calc_reg_comparator_fifth_inp1_14 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_14, QB=>nx34125, D=>nx22531, CLK=>clk);
   ix34129 : nand03 port map ( Y=>nx34128, A0=>label_9_output_14, A1=>
      nx41577, A2=>nx41587);
   labelsregfile_label9_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_9_output_14, QB=>OPEN, D=>nx22521, CLK=>clk, R=>rst);
   lat_label_9_input_14 : latch port map ( Q=>label_9_input_14, D=>nx5512, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_14 : dffr port map ( Q=>
      label_9_input_state_machine_14, QB=>OPEN, D=>nx22251, CLK=>clk, R=>rst
   );
   ix5509 : xnor2 port map ( Y=>nx5508, A0=>nx5504, A1=>nx34755);
   ix5505 : oai22 port map ( Y=>nx5504, A0=>nx34139, A1=>nx34744, B0=>
      nx34754, B1=>nx34513);
   ix34140 : aoi22 port map ( Y=>nx34139, A0=>label_9_output_12, A1=>
      booth_booth_integration_output_8_24, B0=>nx5440, B1=>nx18291);
   labelsregfile_label9_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_9_output_12, QB=>OPEN, D=>nx22491, CLK=>clk, R=>rst);
   lat_label_9_input_12 : latch port map ( Q=>label_9_input_12, D=>nx5454, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_12 : dffr port map ( Q=>
      label_9_input_state_machine_12, QB=>OPEN, D=>nx22481, CLK=>clk, R=>rst
   );
   ix5451 : xnor2 port map ( Y=>nx5450, A0=>nx5440, A1=>nx34740);
   ix5441 : oai22 port map ( Y=>nx5440, A0=>nx34150, A1=>nx34729, B0=>
      nx34739, B1=>nx34477);
   ix34151 : aoi22 port map ( Y=>nx34150, A0=>label_9_output_10, A1=>
      booth_booth_integration_output_8_22, B0=>nx5376, B1=>nx18287);
   labelsregfile_label9_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_9_output_10, QB=>OPEN, D=>nx22451, CLK=>clk, R=>rst);
   lat_label_9_input_10 : latch port map ( Q=>label_9_input_10, D=>nx5390, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_10 : dffr port map ( Q=>
      label_9_input_state_machine_10, QB=>OPEN, D=>nx22441, CLK=>clk, R=>rst
   );
   ix5387 : xnor2 port map ( Y=>nx5386, A0=>nx5376, A1=>nx34725);
   ix5377 : oai22 port map ( Y=>nx5376, A0=>nx34161, A1=>nx34714, B0=>
      nx34724, B1=>nx34441);
   ix34162 : aoi22 port map ( Y=>nx34161, A0=>label_9_output_8, A1=>
      booth_booth_integration_output_8_20, B0=>nx5312, B1=>nx18284);
   labelsregfile_label9_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_9_output_8, QB=>OPEN, D=>nx22411, CLK=>clk, R=>rst);
   lat_label_9_input_8 : latch port map ( Q=>label_9_input_8, D=>nx5326, CLK
      =>nx41671);
   reg_label_9_input_state_machine_8 : dffr port map ( Q=>
      label_9_input_state_machine_8, QB=>OPEN, D=>nx22401, CLK=>clk, R=>rst
   );
   ix5323 : xnor2 port map ( Y=>nx5322, A0=>nx5312, A1=>nx34710);
   ix5313 : oai22 port map ( Y=>nx5312, A0=>nx34172, A1=>nx34699, B0=>
      nx34709, B1=>nx34403);
   ix34173 : aoi22 port map ( Y=>nx34172, A0=>label_9_output_6, A1=>
      booth_booth_integration_output_8_18, B0=>nx5248, B1=>nx18282);
   labelsregfile_label9_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_9_output_6, QB=>OPEN, D=>nx22371, CLK=>clk, R=>rst);
   lat_label_9_input_6 : latch port map ( Q=>label_9_input_6, D=>nx5262, CLK
      =>nx41671);
   reg_label_9_input_state_machine_6 : dffr port map ( Q=>
      label_9_input_state_machine_6, QB=>OPEN, D=>nx22361, CLK=>clk, R=>rst
   );
   ix5259 : xnor2 port map ( Y=>nx5258, A0=>nx5248, A1=>nx34695);
   ix5249 : oai22 port map ( Y=>nx5248, A0=>nx34183, A1=>nx34684, B0=>
      nx34694, B1=>nx34364);
   ix34184 : aoi22 port map ( Y=>nx34183, A0=>label_9_output_4, A1=>
      booth_booth_integration_output_8_16, B0=>nx5184, B1=>nx18280);
   labelsregfile_label9_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_9_output_4, QB=>OPEN, D=>nx22331, CLK=>clk, R=>rst);
   lat_label_9_input_4 : latch port map ( Q=>label_9_input_4, D=>nx5198, CLK
      =>nx41671);
   reg_label_9_input_state_machine_4 : dffr port map ( Q=>
      label_9_input_state_machine_4, QB=>OPEN, D=>nx22321, CLK=>clk, R=>rst
   );
   ix5195 : xnor2 port map ( Y=>nx5194, A0=>nx5184, A1=>nx34680);
   ix5185 : oai22 port map ( Y=>nx5184, A0=>nx34194, A1=>nx34669, B0=>
      nx34679, B1=>nx34647);
   ix34195 : aoi22 port map ( Y=>nx34194, A0=>label_9_output_2, A1=>
      booth_booth_integration_output_8_14, B0=>nx5120, B1=>nx18277);
   labelsregfile_label9_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_9_output_2, QB=>OPEN, D=>nx22291, CLK=>clk, R=>rst);
   lat_label_9_input_2 : latch port map ( Q=>label_9_input_2, D=>nx5134, CLK
      =>nx41669);
   reg_label_9_input_state_machine_2 : dffr port map ( Q=>
      label_9_input_state_machine_2, QB=>OPEN, D=>nx22281, CLK=>clk, R=>rst
   );
   ix5131 : xnor2 port map ( Y=>nx5130, A0=>nx5120, A1=>nx34665);
   ix5121 : oai22 port map ( Y=>nx5120, A0=>nx34205, A1=>nx34654, B0=>
      nx34664, B1=>nx34650);
   ix34206 : nand02 port map ( Y=>nx34205, A0=>label_9_output_0, A1=>
      booth_booth_integration_output_8_12);
   labelsregfile_label9_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_9_output_0, QB=>OPEN, D=>nx21391, CLK=>clk, R=>rst);
   lat_label_9_input_0 : latch port map ( Q=>label_9_input_0, D=>nx3748, CLK
      =>nx41669);
   ix3749 : oai21 port map ( Y=>nx3748, A0=>nx34211, A1=>nx41429, B0=>
      nx34215);
   reg_label_9_input_state_machine_0 : dffr port map ( Q=>
      label_9_input_state_machine_0, QB=>nx34211, D=>nx21381, CLK=>clk, R=>
      rst);
   ix34216 : oai21 port map ( Y=>nx34215, A0=>
      booth_booth_integration_output_8_12, A1=>label_9_output_0, B0=>nx3736
   );
   booth_booth_integrtaion_8_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_12, QB=>OPEN, D=>nx21371, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_13, QB=>nx34650, D=>nx21361, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_14, QB=>OPEN, D=>nx21351, CLK=>clk, R
      =>rst);
   ix34229 : aoi22 port map ( Y=>nx34228, A0=>nx41795, A1=>nx41847, B0=>
      nx3676, B1=>nx3682);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_reg_output_0, QB=>OPEN, 
      D=>nx20871, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_0, QB=>OPEN, D=>nx20857, CLK
      =>clk, S=>nx41483);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_reg_output_9, QB=>OPEN, 
      D=>nx21051, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_9, QB=>OPEN, D=>nx21041, CLK
      =>clk, R=>nx41483);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12912, QB=>OPEN, D=>nx21031, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_8, QB=>OPEN, D=>nx21021, CLK
      =>clk, R=>nx41483);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12913, QB=>OPEN, D=>nx21011, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_7, QB=>OPEN, D=>nx21001, CLK
      =>clk, R=>nx41483);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12914, QB=>OPEN, D=>nx20991, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_6, QB=>OPEN, D=>nx20981, CLK
      =>clk, R=>nx41483);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12915, QB=>OPEN, D=>nx20971, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_5, QB=>OPEN, D=>nx20961, CLK
      =>clk, R=>nx41481);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12916, QB=>OPEN, D=>nx20951, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_4, QB=>OPEN, D=>nx20941, CLK
      =>clk, R=>nx41481);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12917, QB=>OPEN, D=>nx20931, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_3, QB=>OPEN, D=>nx20921, CLK
      =>clk, R=>nx41481);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12918, QB=>OPEN, D=>nx20911, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_2, QB=>OPEN, D=>nx20901, CLK
      =>clk, R=>nx41481);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12919, QB=>OPEN, D=>nx20891, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_1, QB=>OPEN, D=>nx20881, CLK
      =>clk, R=>nx41481);
   ix20852 : nand02 port map ( Y=>nx20851, A0=>nx42933, A1=>nx41833);
   booth_booth_integrtaion_8_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx34275, D=>nx20851, CLK=>clk, S=>nx41481);
   ix3677 : nand02 port map ( Y=>nx3676, A0=>nx34296, A1=>nx34354);
   ix34297 : oai21 port map ( Y=>nx34296, A0=>nx41859, A1=>nx41855, B0=>
      data_in(128));
   ix21182 : oai21 port map ( Y=>nx21181, A0=>nx34301, A1=>nx42497, B0=>
      nx34303);
   booth_booth_integrtaion_8_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx34301, D=>nx21181, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12263, QB=>nx34352, D=>nx21171, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12262, QB=>OPEN, D=>nx21161, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12261, QB=>OPEN, D=>nx21151, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12260, QB=>OPEN, D=>nx21141, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12259, QB=>OPEN, D=>nx21131, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12258, QB=>OPEN, D=>nx21121, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12257, QB=>OPEN, D=>nx21111, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12256, QB=>OPEN, D=>nx21101, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12255, QB=>OPEN, D=>nx21091, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12254, QB=>OPEN, D=>nx21081, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12253, QB=>OPEN, D=>nx21071, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12252, QB=>OPEN, D=>nx21061, CLK=>clk, R=>rst);
   ix34359 : xnor2 port map ( Y=>nx34358, A0=>nx3146, A1=>nx18215);
   ix21322 : oai21 port map ( Y=>nx21321, A0=>nx34364, A1=>nx42497, B0=>
      nx34366);
   booth_booth_integrtaion_8_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_17, QB=>nx34364, D=>nx21321, CLK=>clk, 
      R=>rst);
   ix34367 : nand03 port map ( Y=>nx34366, A0=>nx42505, A1=>nx3654, A2=>
      nx42501);
   ix3655 : xnor2 port map ( Y=>nx3654, A0=>nx34369, A1=>nx18217);
   ix34370 : aoi22 port map ( Y=>nx34369, A0=>
      booth_booth_integration_output_8_17, A1=>nx3170, B0=>nx3146, B1=>
      nx18215);
   ix3161 : nor02_2x port map ( Y=>nx3160, A0=>data_in(128), A1=>
      data_in(129));
   ix21312 : oai21 port map ( Y=>nx21311, A0=>nx34384, A1=>nx42497, B0=>
      nx34386);
   booth_booth_integrtaion_8_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_18, QB=>nx34384, D=>nx21311, CLK=>clk, 
      R=>rst);
   ix34387 : nand03 port map ( Y=>nx34386, A0=>nx42505, A1=>nx3642, A2=>
      nx42501);
   ix3643 : xnor2 port map ( Y=>nx3642, A0=>nx3198, A1=>nx34399);
   ix3199 : oai22 port map ( Y=>nx3198, A0=>nx34369, A1=>nx34390, B0=>
      nx34384, B1=>nx42509);
   ix34393 : aoi32 port map ( Y=>nx34392, A0=>nx3180, A1=>nx41859, A2=>
      nx34395, B0=>data_in(130), B1=>nx41855);
   ix3181 : oai21 port map ( Y=>nx3180, A0=>data_in(128), A1=>data_in(129), 
      B0=>data_in(130));
   ix21302 : oai21 port map ( Y=>nx21301, A0=>nx34403, A1=>nx42497, B0=>
      nx34405);
   booth_booth_integrtaion_8_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_19, QB=>nx34403, D=>nx21301, CLK=>clk, 
      R=>rst);
   ix34406 : nand03 port map ( Y=>nx34405, A0=>nx42505, A1=>nx3630, A2=>
      nx42501);
   ix3631 : xnor2 port map ( Y=>nx3630, A0=>nx34408, A1=>nx18221);
   ix34409 : aoi22 port map ( Y=>nx34408, A0=>
      booth_booth_integration_output_8_19, A1=>nx3218, B0=>nx3198, B1=>
      nx18219);
   ix3219 : oai32 port map ( Y=>nx3218, A0=>nx34411, A1=>nx34374, A2=>nx3208, 
      B0=>nx34414, B1=>nx34379);
   ix3185 : nor03_2x port map ( Y=>nx3184, A0=>data_in(130), A1=>
      data_in(128), A2=>data_in(129));
   ix34415 : inv01 port map ( Y=>nx34414, A=>data_in(131));
   ix3209 : nor04 port map ( Y=>nx3208, A0=>data_in(131), A1=>data_in(130), 
      A2=>data_in(128), A3=>data_in(129));
   ix34423 : xnor2 port map ( Y=>nx34422, A0=>nx3246, A1=>nx18223);
   ix3247 : oai22 port map ( Y=>nx3246, A0=>nx34408, A1=>nx34425, B0=>
      nx34436, B1=>nx42511);
   ix34428 : aoi32 port map ( Y=>nx34427, A0=>nx3228, A1=>nx41859, A2=>
      nx34432, B0=>data_in(132), B1=>nx41855);
   ix3229 : nand02 port map ( Y=>nx3228, A0=>nx34430, A1=>data_in(132));
   ix34433 : nand02 port map ( Y=>nx34432, A0=>nx34434, A1=>nx3208);
   ix34435 : inv01 port map ( Y=>nx34434, A=>data_in(132));
   booth_booth_integrtaion_8_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_20, QB=>nx34436, D=>nx21291, CLK=>clk, 
      R=>rst);
   ix21282 : oai21 port map ( Y=>nx21281, A0=>nx34441, A1=>nx42497, B0=>
      nx34443);
   booth_booth_integrtaion_8_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_21, QB=>nx34441, D=>nx21281, CLK=>clk, 
      R=>rst);
   ix34444 : nand03 port map ( Y=>nx34443, A0=>nx42505, A1=>nx3606, A2=>
      nx42501);
   ix3607 : xnor2 port map ( Y=>nx3606, A0=>nx34446, A1=>nx18225);
   ix34447 : aoi22 port map ( Y=>nx34446, A0=>
      booth_booth_integration_output_8_21, A1=>nx3266, B0=>nx3246, B1=>
      nx18223);
   ix3257 : nor02_2x port map ( Y=>nx3256, A0=>data_in(133), A1=>nx34432);
   ix34459 : xnor2 port map ( Y=>nx34458, A0=>nx3294, A1=>nx18227);
   ix3295 : oai22 port map ( Y=>nx3294, A0=>nx34446, A1=>nx34461, B0=>
      nx34472, B1=>nx42513);
   ix34464 : aoi32 port map ( Y=>nx34463, A0=>nx3276, A1=>nx41859, A2=>
      nx34468, B0=>data_in(134), B1=>nx41855);
   ix3277 : nand02 port map ( Y=>nx3276, A0=>nx34466, A1=>data_in(134));
   ix34469 : nand02 port map ( Y=>nx34468, A0=>nx34470, A1=>nx3256);
   ix34471 : inv01 port map ( Y=>nx34470, A=>data_in(134));
   booth_booth_integrtaion_8_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_22, QB=>nx34472, D=>nx21271, CLK=>clk, 
      R=>rst);
   ix21262 : oai21 port map ( Y=>nx21261, A0=>nx34477, A1=>nx42499, B0=>
      nx34479);
   booth_booth_integrtaion_8_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_23, QB=>nx34477, D=>nx21261, CLK=>clk, 
      R=>rst);
   ix34480 : nand03 port map ( Y=>nx34479, A0=>nx42505, A1=>nx3582, A2=>
      nx42501);
   ix3583 : xnor2 port map ( Y=>nx3582, A0=>nx34482, A1=>nx18228);
   ix34483 : aoi22 port map ( Y=>nx34482, A0=>
      booth_booth_integration_output_8_23, A1=>nx3314, B0=>nx3294, B1=>
      nx18227);
   ix3305 : nor02_2x port map ( Y=>nx3304, A0=>data_in(135), A1=>nx34468);
   ix34495 : xnor2 port map ( Y=>nx34494, A0=>nx3342, A1=>nx18229);
   ix3343 : oai22 port map ( Y=>nx3342, A0=>nx34482, A1=>nx34497, B0=>
      nx34508, B1=>nx42515);
   ix34500 : aoi32 port map ( Y=>nx34499, A0=>nx3324, A1=>nx41859, A2=>
      nx34504, B0=>data_in(136), B1=>nx41855);
   ix3325 : nand02 port map ( Y=>nx3324, A0=>nx34502, A1=>data_in(136));
   ix34505 : nand02 port map ( Y=>nx34504, A0=>nx34506, A1=>nx3304);
   ix34507 : inv01 port map ( Y=>nx34506, A=>data_in(136));
   booth_booth_integrtaion_8_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_24, QB=>nx34508, D=>nx21251, CLK=>clk, 
      R=>rst);
   ix21242 : oai21 port map ( Y=>nx21241, A0=>nx34513, A1=>nx42499, B0=>
      nx34515);
   booth_booth_integrtaion_8_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_25, QB=>nx34513, D=>nx21241, CLK=>clk, 
      R=>rst);
   ix34516 : nand03 port map ( Y=>nx34515, A0=>nx42505, A1=>nx3558, A2=>
      nx42501);
   ix3559 : xnor2 port map ( Y=>nx3558, A0=>nx34518, A1=>nx18230);
   ix34519 : aoi22 port map ( Y=>nx34518, A0=>
      booth_booth_integration_output_8_25, A1=>nx3362, B0=>nx3342, B1=>
      nx18229);
   ix3353 : nor02_2x port map ( Y=>nx3352, A0=>data_in(137), A1=>nx34504);
   ix34531 : xnor2 port map ( Y=>nx34530, A0=>nx3390, A1=>nx18231);
   ix3391 : oai22 port map ( Y=>nx3390, A0=>nx34518, A1=>nx34533, B0=>
      nx34544, B1=>nx42517);
   ix34536 : aoi32 port map ( Y=>nx34535, A0=>nx3372, A1=>nx41859, A2=>
      nx34540, B0=>data_in(138), B1=>nx41855);
   ix3373 : nand02 port map ( Y=>nx3372, A0=>nx34538, A1=>data_in(138));
   ix34541 : nand02 port map ( Y=>nx34540, A0=>nx34542, A1=>nx3352);
   ix34543 : inv01 port map ( Y=>nx34542, A=>data_in(138));
   booth_booth_integrtaion_8_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_26, QB=>nx34544, D=>nx21231, CLK=>clk, 
      R=>rst);
   ix21222 : oai21 port map ( Y=>nx21221, A0=>nx34549, A1=>nx42499, B0=>
      nx34551);
   booth_booth_integrtaion_8_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_27, QB=>nx34549, D=>nx21221, CLK=>clk, 
      R=>rst);
   ix34552 : nand03 port map ( Y=>nx34551, A0=>nx43197, A1=>nx3534, A2=>
      nx42501);
   ix3535 : xnor2 port map ( Y=>nx3534, A0=>nx34554, A1=>nx18232);
   ix34555 : aoi22 port map ( Y=>nx34554, A0=>
      booth_booth_integration_output_8_27, A1=>nx3410, B0=>nx3390, B1=>
      nx18231);
   ix3401 : nor02_2x port map ( Y=>nx3400, A0=>data_in(139), A1=>nx34540);
   ix34567 : xnor2 port map ( Y=>nx34566, A0=>nx3438, A1=>nx18233);
   ix3439 : oai22 port map ( Y=>nx3438, A0=>nx34554, A1=>nx34569, B0=>
      nx34580, B1=>nx42519);
   ix34572 : aoi32 port map ( Y=>nx34571, A0=>nx3420, A1=>nx41861, A2=>
      nx34576, B0=>data_in(140), B1=>nx41855);
   ix3421 : nand02 port map ( Y=>nx3420, A0=>nx34574, A1=>data_in(140));
   ix34577 : nand02 port map ( Y=>nx34576, A0=>nx34578, A1=>nx3400);
   ix34579 : inv01 port map ( Y=>nx34578, A=>data_in(140));
   booth_booth_integrtaion_8_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12251, QB=>nx34580, D=>nx21211, CLK=>clk, R=>rst);
   ix21202 : oai21 port map ( Y=>nx21201, A0=>nx34585, A1=>nx42499, B0=>
      nx34587);
   booth_booth_integrtaion_8_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12250, QB=>nx34585, D=>nx21201, CLK=>clk, R=>rst);
   ix34588 : nand03 port map ( Y=>nx34587, A0=>nx43197, A1=>nx3510, A2=>
      nx42499);
   ix3511 : xnor2 port map ( Y=>nx3510, A0=>nx34590, A1=>nx18235);
   ix34591 : aoi22 port map ( Y=>nx34590, A0=>booth_output_29_dup_12250, A1
      =>nx3458, B0=>nx3438, B1=>nx18233);
   ix3449 : nor02_2x port map ( Y=>nx3448, A0=>data_in(141), A1=>nx34576);
   ix21192 : oai21 port map ( Y=>nx21191, A0=>nx34601, A1=>nx42499, B0=>
      nx34603);
   booth_booth_integrtaion_8_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx34601, D=>nx21191, CLK=>clk, R=>rst);
   ix34604 : nand03 port map ( Y=>nx34603, A0=>nx43197, A1=>nx3498, A2=>
      nx42499);
   ix3499 : xnor2 port map ( Y=>nx3498, A0=>nx3486, A1=>nx34618);
   ix3487 : oai22 port map ( Y=>nx3486, A0=>nx34590, A1=>nx34607, B0=>
      nx34601, B1=>nx42521);
   ix34610 : aoi32 port map ( Y=>nx34609, A0=>nx3468, A1=>nx41861, A2=>
      nx34614, B0=>data_in(142), B1=>nx41857);
   ix3469 : nand02 port map ( Y=>nx3468, A0=>nx34612, A1=>data_in(142));
   ix34615 : nand02 port map ( Y=>nx34614, A0=>nx34616, A1=>nx3448);
   ix34617 : inv01 port map ( Y=>nx34616, A=>data_in(142));
   ix3495 : oai22 port map ( Y=>nx3494, A0=>nx34374, A1=>nx34621, B0=>
      nx34623, B1=>nx34379);
   ix34622 : xnor2 port map ( Y=>nx34621, A0=>data_in(143), A1=>nx34614);
   ix34624 : inv01 port map ( Y=>nx34623, A=>data_in(143));
   ix34626 : aoi32 port map ( Y=>nx34625, A0=>nx3444, A1=>nx41861, A2=>
      nx34612, B0=>data_in(141), B1=>nx41857);
   ix3445 : nand02 port map ( Y=>nx3444, A0=>nx34576, A1=>data_in(141));
   ix34629 : aoi32 port map ( Y=>nx34628, A0=>nx3396, A1=>nx41861, A2=>
      nx34574, B0=>data_in(139), B1=>nx41857);
   ix3397 : nand02 port map ( Y=>nx3396, A0=>nx34540, A1=>data_in(139));
   ix34632 : aoi32 port map ( Y=>nx34631, A0=>nx3348, A1=>nx41861, A2=>
      nx34538, B0=>data_in(137), B1=>nx41857);
   ix3349 : nand02 port map ( Y=>nx3348, A0=>nx34504, A1=>data_in(137));
   ix34635 : aoi32 port map ( Y=>nx34634, A0=>nx3300, A1=>nx41861, A2=>
      nx34502, B0=>data_in(135), B1=>nx41857);
   ix3301 : nand02 port map ( Y=>nx3300, A0=>nx34468, A1=>data_in(135));
   ix34638 : aoi32 port map ( Y=>nx34637, A0=>nx3252, A1=>nx41863, A2=>
      nx34466, B0=>data_in(133), B1=>nx41857);
   ix3253 : nand02 port map ( Y=>nx3252, A0=>nx34432, A1=>data_in(133));
   ix34641 : aoi32 port map ( Y=>nx34640, A0=>nx3154, A1=>nx41863, A2=>
      nx34643, B0=>data_in(129), B1=>nx41857);
   ix3155 : nand02 port map ( Y=>nx3154, A0=>data_in(129), A1=>data_in(128)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_16, QB=>nx34354, D=>nx21331, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_15, QB=>nx34647, D=>nx21341, CLK=>clk, 
      R=>rst);
   ix3737 : aoi21 port map ( Y=>nx3736, A0=>label_9_output_0, A1=>
      booth_booth_integration_output_8_12, B0=>nx43519);
   labelsregfile_label9_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_9_output_1, QB=>nx34664, D=>nx22271, CLK=>clk, R=>rst);
   lat_label_9_input_1 : latch port map ( Q=>label_9_input_1, D=>nx5102, CLK
      =>nx41669);
   reg_label_9_input_state_machine_1 : dffr port map ( Q=>
      label_9_input_state_machine_1, QB=>OPEN, D=>nx22261, CLK=>clk, R=>rst
   );
   ix5099 : xor2 port map ( Y=>nx5098, A0=>nx34205, A1=>nx34654);
   ix34666 : xnor2 port map ( Y=>nx34665, A0=>
      booth_booth_integration_output_8_14, A1=>label_9_output_2);
   labelsregfile_label9_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_9_output_3, QB=>nx34679, D=>nx22311, CLK=>clk, R=>rst);
   lat_label_9_input_3 : latch port map ( Q=>label_9_input_3, D=>nx5166, CLK
      =>nx41671);
   reg_label_9_input_state_machine_3 : dffr port map ( Q=>
      label_9_input_state_machine_3, QB=>OPEN, D=>nx22301, CLK=>clk, R=>rst
   );
   ix5163 : xor2 port map ( Y=>nx5162, A0=>nx34194, A1=>nx34669);
   labelsregfile_label9_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_9_output_5, QB=>nx34694, D=>nx22351, CLK=>clk, R=>rst);
   lat_label_9_input_5 : latch port map ( Q=>label_9_input_5, D=>nx5230, CLK
      =>nx41671);
   reg_label_9_input_state_machine_5 : dffr port map ( Q=>
      label_9_input_state_machine_5, QB=>OPEN, D=>nx22341, CLK=>clk, R=>rst
   );
   ix5227 : xor2 port map ( Y=>nx5226, A0=>nx34183, A1=>nx34684);
   labelsregfile_label9_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_9_output_7, QB=>nx34709, D=>nx22391, CLK=>clk, R=>rst);
   lat_label_9_input_7 : latch port map ( Q=>label_9_input_7, D=>nx5294, CLK
      =>nx41671);
   reg_label_9_input_state_machine_7 : dffr port map ( Q=>
      label_9_input_state_machine_7, QB=>OPEN, D=>nx22381, CLK=>clk, R=>rst
   );
   ix5291 : xor2 port map ( Y=>nx5290, A0=>nx34172, A1=>nx34699);
   labelsregfile_label9_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_9_output_9, QB=>nx34724, D=>nx22431, CLK=>clk, R=>rst);
   lat_label_9_input_9 : latch port map ( Q=>label_9_input_9, D=>nx5358, CLK
      =>nx41671);
   reg_label_9_input_state_machine_9 : dffr port map ( Q=>
      label_9_input_state_machine_9, QB=>OPEN, D=>nx22421, CLK=>clk, R=>rst
   );
   ix5355 : xor2 port map ( Y=>nx5354, A0=>nx34161, A1=>nx34714);
   labelsregfile_label9_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_9_output_11, QB=>nx34739, D=>nx22471, CLK=>clk, R=>rst);
   lat_label_9_input_11 : latch port map ( Q=>label_9_input_11, D=>nx5422, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_11 : dffr port map ( Q=>
      label_9_input_state_machine_11, QB=>OPEN, D=>nx22461, CLK=>clk, R=>rst
   );
   ix5419 : xor2 port map ( Y=>nx5418, A0=>nx34150, A1=>nx34729);
   labelsregfile_label9_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_9_output_13, QB=>nx34754, D=>nx22511, CLK=>clk, R=>rst);
   lat_label_9_input_13 : latch port map ( Q=>label_9_input_13, D=>nx5486, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_13 : dffr port map ( Q=>
      label_9_input_state_machine_13, QB=>OPEN, D=>nx22501, CLK=>clk, R=>rst
   );
   ix5483 : xor2 port map ( Y=>nx5482, A0=>nx34139, A1=>nx34744);
   ix22242 : oai21 port map ( Y=>nx22241, A0=>nx34760, A1=>nx41587, B0=>
      nx34762);
   max_calc_reg_comparator_fifth_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx34760, D=>nx22241, CLK=>clk);
   ix34763 : nand03 port map ( Y=>nx34762, A0=>label_10_output_14, A1=>
      nx41577, A2=>nx41587);
   ix5979 : xnor2 port map ( Y=>nx5978, A0=>nx34765, A1=>nx5976);
   ix34766 : aoi22 port map ( Y=>nx34765, A0=>nx34760, A1=>
      max_calc_comparator_fifth_inp1_14, B0=>nx5532, B1=>nx5886);
   ix5887 : oai22 port map ( Y=>nx5886, A0=>nx34769, A1=>nx34782, B0=>
      max_calc_comparator_fifth_inp2_13, B1=>nx34777);
   ix22542 : oai21 port map ( Y=>nx22541, A0=>nx34773, A1=>nx41587, B0=>
      nx34775);
   max_calc_reg_comparator_fifth_inp2_13 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_13, QB=>nx34773, D=>nx22541, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_13 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_13, QB=>nx34777, D=>nx22551, CLK=>clk);
   ix22552 : oai21 port map ( Y=>nx22551, A0=>nx34777, A1=>nx41587, B0=>
      nx34780);
   ix34783 : aoi22 port map ( Y=>nx34782, A0=>nx34784, A1=>
      max_calc_comparator_fifth_inp1_12, B0=>nx5568, B1=>nx5870);
   max_calc_reg_comparator_fifth_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx34784, D=>nx22561, CLK=>clk);
   ix22562 : oai21 port map ( Y=>nx22561, A0=>nx34784, A1=>nx41589, B0=>
      nx34787);
   ix34788 : nand03 port map ( Y=>nx34787, A0=>label_10_output_12, A1=>
      nx41577, A2=>nx41589);
   ix22572 : oai21 port map ( Y=>nx22571, A0=>nx34791, A1=>nx41589, B0=>
      nx34793);
   max_calc_reg_comparator_fifth_inp1_12 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_12, QB=>nx34791, D=>nx22571, CLK=>clk);
   ix34794 : nand03 port map ( Y=>nx34793, A0=>label_9_output_12, A1=>
      nx41577, A2=>nx41589);
   ix5871 : oai22 port map ( Y=>nx5870, A0=>nx34797, A1=>nx34810, B0=>
      max_calc_comparator_fifth_inp2_11, B1=>nx34805);
   ix22582 : oai21 port map ( Y=>nx22581, A0=>nx34801, A1=>nx41589, B0=>
      nx34803);
   max_calc_reg_comparator_fifth_inp2_11 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_11, QB=>nx34801, D=>nx22581, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_11 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_11, QB=>nx34805, D=>nx22591, CLK=>clk);
   ix22592 : oai21 port map ( Y=>nx22591, A0=>nx34805, A1=>nx41591, B0=>
      nx34808);
   ix34811 : aoi22 port map ( Y=>nx34810, A0=>nx34812, A1=>
      max_calc_comparator_fifth_inp1_10, B0=>nx5604, B1=>nx5854);
   max_calc_reg_comparator_fifth_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx34812, D=>nx22601, CLK=>clk);
   ix22602 : oai21 port map ( Y=>nx22601, A0=>nx34812, A1=>nx41591, B0=>
      nx34815);
   ix34816 : nand03 port map ( Y=>nx34815, A0=>label_10_output_10, A1=>
      nx41579, A2=>nx41591);
   ix22612 : oai21 port map ( Y=>nx22611, A0=>nx34819, A1=>nx41591, B0=>
      nx34821);
   max_calc_reg_comparator_fifth_inp1_10 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_10, QB=>nx34819, D=>nx22611, CLK=>clk);
   ix34822 : nand03 port map ( Y=>nx34821, A0=>label_9_output_10, A1=>
      nx41579, A2=>nx41591);
   ix5855 : oai22 port map ( Y=>nx5854, A0=>nx34825, A1=>nx34838, B0=>
      max_calc_comparator_fifth_inp2_9, B1=>nx34833);
   ix22622 : oai21 port map ( Y=>nx22621, A0=>nx34829, A1=>nx41591, B0=>
      nx34831);
   max_calc_reg_comparator_fifth_inp2_9 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_9, QB=>nx34829, D=>nx22621, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_9 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_9, QB=>nx34833, D=>nx22631, CLK=>clk);
   ix22632 : oai21 port map ( Y=>nx22631, A0=>nx34833, A1=>nx41593, B0=>
      nx34836);
   ix34839 : aoi22 port map ( Y=>nx34838, A0=>nx34840, A1=>
      max_calc_comparator_fifth_inp1_8, B0=>nx5640, B1=>nx5838);
   max_calc_reg_comparator_fifth_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx34840, D=>nx22641, CLK=>clk);
   ix22642 : oai21 port map ( Y=>nx22641, A0=>nx34840, A1=>nx41593, B0=>
      nx34843);
   ix34844 : nand03 port map ( Y=>nx34843, A0=>label_10_output_8, A1=>
      nx41579, A2=>nx41593);
   ix22652 : oai21 port map ( Y=>nx22651, A0=>nx34847, A1=>nx41593, B0=>
      nx34849);
   max_calc_reg_comparator_fifth_inp1_8 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_8, QB=>nx34847, D=>nx22651, CLK=>clk);
   ix34850 : nand03 port map ( Y=>nx34849, A0=>label_9_output_8, A1=>nx41581, 
      A2=>nx41593);
   ix5839 : oai22 port map ( Y=>nx5838, A0=>nx34853, A1=>nx34866, B0=>
      max_calc_comparator_fifth_inp2_7, B1=>nx34861);
   ix22662 : oai21 port map ( Y=>nx22661, A0=>nx34857, A1=>nx41595, B0=>
      nx34859);
   max_calc_reg_comparator_fifth_inp2_7 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_7, QB=>nx34857, D=>nx22661, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_7 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_7, QB=>nx34861, D=>nx22671, CLK=>clk);
   ix22672 : oai21 port map ( Y=>nx22671, A0=>nx34861, A1=>nx41595, B0=>
      nx34864);
   ix34867 : aoi22 port map ( Y=>nx34866, A0=>nx34868, A1=>
      max_calc_comparator_fifth_inp1_6, B0=>nx5676, B1=>nx5822);
   max_calc_reg_comparator_fifth_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx34868, D=>nx22681, CLK=>clk);
   ix22682 : oai21 port map ( Y=>nx22681, A0=>nx34868, A1=>nx41595, B0=>
      nx34871);
   ix34872 : nand03 port map ( Y=>nx34871, A0=>label_10_output_6, A1=>
      nx41581, A2=>nx41595);
   ix22692 : oai21 port map ( Y=>nx22691, A0=>nx34875, A1=>nx41595, B0=>
      nx34877);
   max_calc_reg_comparator_fifth_inp1_6 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_6, QB=>nx34875, D=>nx22691, CLK=>clk);
   ix34878 : nand03 port map ( Y=>nx34877, A0=>label_9_output_6, A1=>nx41581, 
      A2=>nx41597);
   ix5823 : oai22 port map ( Y=>nx5822, A0=>nx34881, A1=>nx34894, B0=>
      max_calc_comparator_fifth_inp2_5, B1=>nx34889);
   ix22702 : oai21 port map ( Y=>nx22701, A0=>nx34885, A1=>nx41597, B0=>
      nx34887);
   max_calc_reg_comparator_fifth_inp2_5 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_5, QB=>nx34885, D=>nx22701, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_5 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_5, QB=>nx34889, D=>nx22711, CLK=>clk);
   ix22712 : oai21 port map ( Y=>nx22711, A0=>nx34889, A1=>nx41597, B0=>
      nx34892);
   ix34895 : aoi22 port map ( Y=>nx34894, A0=>nx34896, A1=>
      max_calc_comparator_fifth_inp1_4, B0=>nx5712, B1=>nx5806);
   max_calc_reg_comparator_fifth_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx34896, D=>nx22721, CLK=>clk);
   ix22722 : oai21 port map ( Y=>nx22721, A0=>nx34896, A1=>nx41597, B0=>
      nx34899);
   ix34900 : nand03 port map ( Y=>nx34899, A0=>label_10_output_4, A1=>
      nx41583, A2=>nx41597);
   ix22732 : oai21 port map ( Y=>nx22731, A0=>nx34903, A1=>nx41599, B0=>
      nx34905);
   max_calc_reg_comparator_fifth_inp1_4 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_4, QB=>nx34903, D=>nx22731, CLK=>clk);
   ix34906 : nand03 port map ( Y=>nx34905, A0=>label_9_output_4, A1=>nx41583, 
      A2=>nx41599);
   ix5807 : oai22 port map ( Y=>nx5806, A0=>nx34909, A1=>nx34922, B0=>
      max_calc_comparator_fifth_inp2_3, B1=>nx34917);
   ix22742 : oai21 port map ( Y=>nx22741, A0=>nx34913, A1=>nx41599, B0=>
      nx34915);
   max_calc_reg_comparator_fifth_inp2_3 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_3, QB=>nx34913, D=>nx22741, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_3 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_3, QB=>nx34917, D=>nx22751, CLK=>clk);
   ix22752 : oai21 port map ( Y=>nx22751, A0=>nx34917, A1=>nx41599, B0=>
      nx34920);
   ix34923 : aoi22 port map ( Y=>nx34922, A0=>nx34924, A1=>
      max_calc_comparator_fifth_inp1_2, B0=>nx5748, B1=>nx5790);
   max_calc_reg_comparator_fifth_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx34924, D=>nx22761, CLK=>clk);
   ix22762 : oai21 port map ( Y=>nx22761, A0=>nx34924, A1=>nx41599, B0=>
      nx34927);
   ix34928 : nand03 port map ( Y=>nx34927, A0=>label_10_output_2, A1=>
      nx41583, A2=>nx41601);
   ix22772 : oai21 port map ( Y=>nx22771, A0=>nx34931, A1=>nx41601, B0=>
      nx34933);
   max_calc_reg_comparator_fifth_inp1_2 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_2, QB=>nx34931, D=>nx22771, CLK=>clk);
   ix34934 : nand03 port map ( Y=>nx34933, A0=>label_9_output_2, A1=>nx41583, 
      A2=>nx41601);
   ix5791 : oai21 port map ( Y=>nx5790, A0=>max_calc_comparator_fifth_inp2_1, 
      A1=>nx34943, B0=>nx34948);
   ix22782 : oai21 port map ( Y=>nx22781, A0=>nx34939, A1=>nx41601, B0=>
      nx34941);
   max_calc_reg_comparator_fifth_inp2_1 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_1, QB=>nx34939, D=>nx22781, CLK=>clk);
   max_calc_reg_comparator_fifth_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx34943, D=>nx22791, CLK=>clk);
   ix22792 : oai21 port map ( Y=>nx22791, A0=>nx34943, A1=>nx41601, B0=>
      nx34946);
   ix34949 : oai21 port map ( Y=>nx34948, A0=>nx34950, A1=>
      max_calc_comparator_fifth_inp1_0, B0=>nx5766);
   max_calc_reg_comparator_fifth_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx34950, D=>nx22801, CLK=>clk);
   ix22802 : oai21 port map ( Y=>nx22801, A0=>nx34950, A1=>nx41603, B0=>
      nx34953);
   ix34954 : nand03 port map ( Y=>nx34953, A0=>label_10_output_0, A1=>
      nx41585, A2=>nx41603);
   ix21402 : oai21 port map ( Y=>nx21401, A0=>nx34957, A1=>nx41603, B0=>
      nx34959);
   max_calc_reg_comparator_fifth_inp1_0 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_0, QB=>nx34957, D=>nx21401, CLK=>clk);
   ix34960 : nand03 port map ( Y=>nx34959, A0=>label_9_output_0, A1=>nx41585, 
      A2=>nx41603);
   ix22832 : oai21 port map ( Y=>nx22831, A0=>nx34965, A1=>nx41603, B0=>
      nx34967);
   max_calc_reg_comparator_fifth_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx34965, D=>nx22831, CLK=>clk);
   ix22862 : oai21 port map ( Y=>nx22861, A0=>nx34971, A1=>nx41603, B0=>
      nx34973);
   max_calc_reg_comparator_fifth_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx34971, D=>nx22861, CLK=>clk);
   lat_label_9_input_15 : latch port map ( Q=>label_9_input_15, D=>nx5956, 
      CLK=>nx41673);
   reg_label_9_input_state_machine_15 : dffr port map ( Q=>
      label_9_input_state_machine_15, QB=>OPEN, D=>nx22841, CLK=>clk, R=>rst
   );
   ix5953 : xnor2 port map ( Y=>nx5952, A0=>nx34983, A1=>nx5950);
   ix34984 : aoi22 port map ( Y=>nx34983, A0=>label_9_output_14, A1=>
      booth_booth_integration_output_8_26, B0=>nx5504, B1=>nx5506);
   labelsregfile_label9_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_9_output_15, QB=>nx34987, D=>nx22851, CLK=>clk, R=>rst);
   ix34994 : nand04 port map ( Y=>nx34993, A0=>nx31955, A1=>max_calc_start, 
      A2=>nx42925, A3=>max_calc_state_0);
   max_calc_reg_comparator_first_inp2_14 : dff port map ( Q=>
      max_calc_comparator_first_inp2_14, QB=>nx40326, D=>nx30451, CLK=>clk);
   labelsregfile_label2_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_2_output_14, QB=>OPEN, D=>nx23711, CLK=>clk, R=>rst);
   lat_label_2_input_14 : latch port map ( Q=>label_2_input_14, D=>nx7302, 
      CLK=>nx41677);
   reg_label_2_input_state_machine_14 : dffr port map ( Q=>
      label_2_input_state_machine_14, QB=>OPEN, D=>nx22891, CLK=>clk, R=>rst
   );
   ix7299 : xnor2 port map ( Y=>nx7298, A0=>nx7294, A1=>nx35625);
   ix7295 : oai22 port map ( Y=>nx7294, A0=>nx35009, A1=>nx35614, B0=>
      nx35624, B1=>nx35383);
   ix35010 : aoi22 port map ( Y=>nx35009, A0=>label_2_output_12, A1=>
      booth_booth_integration_output_1_24, B0=>nx7230, B1=>nx18334);
   labelsregfile_label2_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_2_output_12, QB=>OPEN, D=>nx23681, CLK=>clk, R=>rst);
   lat_label_2_input_12 : latch port map ( Q=>label_2_input_12, D=>nx7244, 
      CLK=>nx41677);
   reg_label_2_input_state_machine_12 : dffr port map ( Q=>
      label_2_input_state_machine_12, QB=>OPEN, D=>nx23671, CLK=>clk, R=>rst
   );
   ix7241 : xnor2 port map ( Y=>nx7240, A0=>nx7230, A1=>nx35610);
   ix7231 : oai22 port map ( Y=>nx7230, A0=>nx35020, A1=>nx35599, B0=>
      nx35609, B1=>nx35347);
   ix35021 : aoi22 port map ( Y=>nx35020, A0=>label_2_output_10, A1=>
      booth_booth_integration_output_1_22, B0=>nx7166, B1=>nx18332);
   labelsregfile_label2_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_2_output_10, QB=>OPEN, D=>nx23641, CLK=>clk, R=>rst);
   lat_label_2_input_10 : latch port map ( Q=>label_2_input_10, D=>nx7180, 
      CLK=>nx41677);
   reg_label_2_input_state_machine_10 : dffr port map ( Q=>
      label_2_input_state_machine_10, QB=>OPEN, D=>nx23631, CLK=>clk, R=>rst
   );
   ix7177 : xnor2 port map ( Y=>nx7176, A0=>nx7166, A1=>nx35595);
   ix7167 : oai22 port map ( Y=>nx7166, A0=>nx35031, A1=>nx35584, B0=>
      nx35594, B1=>nx35311);
   ix35032 : aoi22 port map ( Y=>nx35031, A0=>label_2_output_8, A1=>
      booth_booth_integration_output_1_20, B0=>nx7102, B1=>nx18329);
   labelsregfile_label2_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_2_output_8, QB=>OPEN, D=>nx23601, CLK=>clk, R=>rst);
   lat_label_2_input_8 : latch port map ( Q=>label_2_input_8, D=>nx7116, CLK
      =>nx41677);
   reg_label_2_input_state_machine_8 : dffr port map ( Q=>
      label_2_input_state_machine_8, QB=>OPEN, D=>nx23591, CLK=>clk, R=>rst
   );
   ix7113 : xnor2 port map ( Y=>nx7112, A0=>nx7102, A1=>nx35580);
   ix7103 : oai22 port map ( Y=>nx7102, A0=>nx35042, A1=>nx35569, B0=>
      nx35579, B1=>nx35273);
   ix35043 : aoi22 port map ( Y=>nx35042, A0=>label_2_output_6, A1=>
      booth_booth_integration_output_1_18, B0=>nx7038, B1=>nx18325);
   labelsregfile_label2_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_2_output_6, QB=>OPEN, D=>nx23561, CLK=>clk, R=>rst);
   lat_label_2_input_6 : latch port map ( Q=>label_2_input_6, D=>nx7052, CLK
      =>nx41675);
   reg_label_2_input_state_machine_6 : dffr port map ( Q=>
      label_2_input_state_machine_6, QB=>OPEN, D=>nx23551, CLK=>clk, R=>rst
   );
   ix7049 : xnor2 port map ( Y=>nx7048, A0=>nx7038, A1=>nx35565);
   ix7039 : oai22 port map ( Y=>nx7038, A0=>nx35053, A1=>nx35554, B0=>
      nx35564, B1=>nx35234);
   ix35054 : aoi22 port map ( Y=>nx35053, A0=>label_2_output_4, A1=>
      booth_booth_integration_output_1_16, B0=>nx6974, B1=>nx18322);
   labelsregfile_label2_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_2_output_4, QB=>OPEN, D=>nx23521, CLK=>clk, R=>rst);
   lat_label_2_input_4 : latch port map ( Q=>label_2_input_4, D=>nx6988, CLK
      =>nx41675);
   reg_label_2_input_state_machine_4 : dffr port map ( Q=>
      label_2_input_state_machine_4, QB=>OPEN, D=>nx23511, CLK=>clk, R=>rst
   );
   ix6985 : xnor2 port map ( Y=>nx6984, A0=>nx6974, A1=>nx35550);
   ix6975 : oai22 port map ( Y=>nx6974, A0=>nx35064, A1=>nx35539, B0=>
      nx35549, B1=>nx35517);
   ix35065 : aoi22 port map ( Y=>nx35064, A0=>label_2_output_2, A1=>
      booth_booth_integration_output_1_14, B0=>nx6910, B1=>nx18320);
   labelsregfile_label2_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_2_output_2, QB=>OPEN, D=>nx23481, CLK=>clk, R=>rst);
   lat_label_2_input_2 : latch port map ( Q=>label_2_input_2, D=>nx6924, CLK
      =>nx41675);
   reg_label_2_input_state_machine_2 : dffr port map ( Q=>
      label_2_input_state_machine_2, QB=>OPEN, D=>nx23471, CLK=>clk, R=>rst
   );
   ix6921 : xnor2 port map ( Y=>nx6920, A0=>nx6910, A1=>nx35535);
   ix6911 : oai22 port map ( Y=>nx6910, A0=>nx35075, A1=>nx35524, B0=>
      nx35534, B1=>nx35520);
   ix35076 : nand02 port map ( Y=>nx35075, A0=>label_2_output_0, A1=>
      booth_booth_integration_output_1_12);
   labelsregfile_label2_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_2_output_0, QB=>OPEN, D=>nx23441, CLK=>clk, R=>rst);
   lat_label_2_input_0 : latch port map ( Q=>label_2_input_0, D=>nx6866, CLK
      =>nx41673);
   ix6867 : oai21 port map ( Y=>nx6866, A0=>nx35081, A1=>nx41435, B0=>
      nx35085);
   reg_label_2_input_state_machine_0 : dffr port map ( Q=>
      label_2_input_state_machine_0, QB=>nx35081, D=>nx23431, CLK=>clk, R=>
      rst);
   ix35086 : oai21 port map ( Y=>nx35085, A0=>
      booth_booth_integration_output_1_12, A1=>label_2_output_0, B0=>nx6854
   );
   booth_booth_integrtaion_1_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_12, QB=>OPEN, D=>nx23421, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_13, QB=>nx35520, D=>nx23411, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_14, QB=>OPEN, D=>nx23401, CLK=>clk, R
      =>rst);
   ix35099 : aoi22 port map ( Y=>nx35098, A0=>nx41795, A1=>nx41919, B0=>
      nx6796, B1=>nx6802);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_reg_output_0, QB=>OPEN, 
      D=>nx22921, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_0, QB=>OPEN, D=>nx22907, CLK
      =>clk, S=>nx41487);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_reg_output_9, QB=>OPEN, 
      D=>nx23101, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_9, QB=>OPEN, D=>nx23091, CLK
      =>clk, R=>nx41487);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12716, QB=>OPEN, D=>nx23081, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_8, QB=>OPEN, D=>nx23071, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12717, QB=>OPEN, D=>nx23061, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_7, QB=>OPEN, D=>nx23051, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12718, QB=>OPEN, D=>nx23041, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_6, QB=>OPEN, D=>nx23031, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12719, QB=>OPEN, D=>nx23021, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_5, QB=>OPEN, D=>nx23011, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12720, QB=>OPEN, D=>nx23001, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_4, QB=>OPEN, D=>nx22991, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12721, QB=>OPEN, D=>nx22981, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_3, QB=>OPEN, D=>nx22971, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12722, QB=>OPEN, D=>nx22961, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_2, QB=>OPEN, D=>nx22951, CLK
      =>clk, R=>nx41485);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12723, QB=>OPEN, D=>nx22941, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_1, QB=>OPEN, D=>nx22931, CLK
      =>clk, R=>nx41483);
   ix22902 : nand02 port map ( Y=>nx22901, A0=>nx42937, A1=>nx41905);
   booth_booth_integrtaion_1_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx35145, D=>nx22901, CLK=>clk, S=>nx41483);
   ix6797 : nand02 port map ( Y=>nx6796, A0=>nx35166, A1=>nx35224);
   ix35167 : oai21 port map ( Y=>nx35166, A0=>nx41931, A1=>nx41927, B0=>
      data_in(16));
   ix23232 : oai21 port map ( Y=>nx23231, A0=>nx35171, A1=>nx42551, B0=>
      nx35173);
   booth_booth_integrtaion_1_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx35171, D=>nx23231, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12130, QB=>nx35222, D=>nx23221, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12129, QB=>OPEN, D=>nx23211, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12128, QB=>OPEN, D=>nx23201, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12127, QB=>OPEN, D=>nx23191, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12126, QB=>OPEN, D=>nx23181, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12125, QB=>OPEN, D=>nx23171, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12124, QB=>OPEN, D=>nx23161, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12123, QB=>OPEN, D=>nx23151, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12122, QB=>OPEN, D=>nx23141, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12121, QB=>OPEN, D=>nx23131, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12120, QB=>OPEN, D=>nx23121, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12119, QB=>OPEN, D=>nx23111, CLK=>clk, R=>rst);
   ix35229 : xnor2 port map ( Y=>nx35228, A0=>nx6266, A1=>nx18297);
   ix23372 : oai21 port map ( Y=>nx23371, A0=>nx35234, A1=>nx42551, B0=>
      nx35236);
   booth_booth_integrtaion_1_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_17, QB=>nx35234, D=>nx23371, CLK=>clk, 
      R=>rst);
   ix35237 : nand03 port map ( Y=>nx35236, A0=>nx42559, A1=>nx6774, A2=>
      nx42555);
   ix6775 : xnor2 port map ( Y=>nx6774, A0=>nx35239, A1=>nx18299);
   ix35240 : aoi22 port map ( Y=>nx35239, A0=>
      booth_booth_integration_output_1_17, A1=>nx6290, B0=>nx6266, B1=>
      nx18297);
   ix6281 : nor02_2x port map ( Y=>nx6280, A0=>data_in(16), A1=>data_in(17)
   );
   ix23362 : oai21 port map ( Y=>nx23361, A0=>nx35254, A1=>nx42551, B0=>
      nx35256);
   booth_booth_integrtaion_1_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_18, QB=>nx35254, D=>nx23361, CLK=>clk, 
      R=>rst);
   ix35257 : nand03 port map ( Y=>nx35256, A0=>nx42559, A1=>nx6762, A2=>
      nx42555);
   ix6763 : xnor2 port map ( Y=>nx6762, A0=>nx6318, A1=>nx35269);
   ix6319 : oai22 port map ( Y=>nx6318, A0=>nx35239, A1=>nx35260, B0=>
      nx35254, B1=>nx42563);
   ix35263 : aoi32 port map ( Y=>nx35262, A0=>nx6300, A1=>nx41931, A2=>
      nx35265, B0=>data_in(18), B1=>nx41927);
   ix6301 : oai21 port map ( Y=>nx6300, A0=>data_in(16), A1=>data_in(17), B0
      =>data_in(18));
   ix23352 : oai21 port map ( Y=>nx23351, A0=>nx35273, A1=>nx42551, B0=>
      nx35275);
   booth_booth_integrtaion_1_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_19, QB=>nx35273, D=>nx23351, CLK=>clk, 
      R=>rst);
   ix35276 : nand03 port map ( Y=>nx35275, A0=>nx42559, A1=>nx6750, A2=>
      nx42555);
   ix6751 : xnor2 port map ( Y=>nx6750, A0=>nx35278, A1=>nx18301);
   ix35279 : aoi22 port map ( Y=>nx35278, A0=>
      booth_booth_integration_output_1_19, A1=>nx6338, B0=>nx6318, B1=>
      nx18300);
   ix6339 : oai32 port map ( Y=>nx6338, A0=>nx35281, A1=>nx35244, A2=>nx6328, 
      B0=>nx35284, B1=>nx35249);
   ix6305 : nor03_2x port map ( Y=>nx6304, A0=>data_in(18), A1=>data_in(16), 
      A2=>data_in(17));
   ix35285 : inv01 port map ( Y=>nx35284, A=>data_in(19));
   ix6329 : nor04 port map ( Y=>nx6328, A0=>data_in(19), A1=>data_in(18), A2
      =>data_in(16), A3=>data_in(17));
   ix35293 : xnor2 port map ( Y=>nx35292, A0=>nx6366, A1=>nx18302);
   ix6367 : oai22 port map ( Y=>nx6366, A0=>nx35278, A1=>nx35295, B0=>
      nx35306, B1=>nx42565);
   ix35298 : aoi32 port map ( Y=>nx35297, A0=>nx6348, A1=>nx41931, A2=>
      nx35302, B0=>data_in(20), B1=>nx41927);
   ix6349 : nand02 port map ( Y=>nx6348, A0=>nx35300, A1=>data_in(20));
   ix35303 : nand02 port map ( Y=>nx35302, A0=>nx35304, A1=>nx6328);
   ix35305 : inv01 port map ( Y=>nx35304, A=>data_in(20));
   booth_booth_integrtaion_1_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_20, QB=>nx35306, D=>nx23341, CLK=>clk, 
      R=>rst);
   ix23332 : oai21 port map ( Y=>nx23331, A0=>nx35311, A1=>nx42551, B0=>
      nx35313);
   booth_booth_integrtaion_1_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_21, QB=>nx35311, D=>nx23331, CLK=>clk, 
      R=>rst);
   ix35314 : nand03 port map ( Y=>nx35313, A0=>nx42559, A1=>nx6726, A2=>
      nx42555);
   ix6727 : xnor2 port map ( Y=>nx6726, A0=>nx35316, A1=>nx18303);
   ix35317 : aoi22 port map ( Y=>nx35316, A0=>
      booth_booth_integration_output_1_21, A1=>nx6386, B0=>nx6366, B1=>
      nx18302);
   ix6377 : nor02_2x port map ( Y=>nx6376, A0=>data_in(21), A1=>nx35302);
   ix35329 : xnor2 port map ( Y=>nx35328, A0=>nx6414, A1=>nx18304);
   ix6415 : oai22 port map ( Y=>nx6414, A0=>nx35316, A1=>nx35331, B0=>
      nx35342, B1=>nx42567);
   ix35334 : aoi32 port map ( Y=>nx35333, A0=>nx6396, A1=>nx41931, A2=>
      nx35338, B0=>data_in(22), B1=>nx41927);
   ix6397 : nand02 port map ( Y=>nx6396, A0=>nx35336, A1=>data_in(22));
   ix35339 : nand02 port map ( Y=>nx35338, A0=>nx35340, A1=>nx6376);
   ix35341 : inv01 port map ( Y=>nx35340, A=>data_in(22));
   booth_booth_integrtaion_1_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_22, QB=>nx35342, D=>nx23321, CLK=>clk, 
      R=>rst);
   ix23312 : oai21 port map ( Y=>nx23311, A0=>nx35347, A1=>nx42553, B0=>
      nx35349);
   booth_booth_integrtaion_1_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_23, QB=>nx35347, D=>nx23311, CLK=>clk, 
      R=>rst);
   ix35350 : nand03 port map ( Y=>nx35349, A0=>nx42559, A1=>nx6702, A2=>
      nx42555);
   ix6703 : xnor2 port map ( Y=>nx6702, A0=>nx35352, A1=>nx18305);
   ix35353 : aoi22 port map ( Y=>nx35352, A0=>
      booth_booth_integration_output_1_23, A1=>nx6434, B0=>nx6414, B1=>
      nx18304);
   ix6425 : nor02_2x port map ( Y=>nx6424, A0=>data_in(23), A1=>nx35338);
   ix35365 : xnor2 port map ( Y=>nx35364, A0=>nx6462, A1=>nx18307);
   ix6463 : oai22 port map ( Y=>nx6462, A0=>nx35352, A1=>nx35367, B0=>
      nx35378, B1=>nx42569);
   ix35370 : aoi32 port map ( Y=>nx35369, A0=>nx6444, A1=>nx41931, A2=>
      nx35374, B0=>data_in(24), B1=>nx41927);
   ix6445 : nand02 port map ( Y=>nx6444, A0=>nx35372, A1=>data_in(24));
   ix35375 : nand02 port map ( Y=>nx35374, A0=>nx35376, A1=>nx6424);
   ix35377 : inv01 port map ( Y=>nx35376, A=>data_in(24));
   booth_booth_integrtaion_1_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_24, QB=>nx35378, D=>nx23301, CLK=>clk, 
      R=>rst);
   ix23292 : oai21 port map ( Y=>nx23291, A0=>nx35383, A1=>nx42553, B0=>
      nx35385);
   booth_booth_integrtaion_1_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_25, QB=>nx35383, D=>nx23291, CLK=>clk, 
      R=>rst);
   ix35386 : nand03 port map ( Y=>nx35385, A0=>nx42559, A1=>nx6678, A2=>
      nx42555);
   ix6679 : xnor2 port map ( Y=>nx6678, A0=>nx35388, A1=>nx18309);
   ix35389 : aoi22 port map ( Y=>nx35388, A0=>
      booth_booth_integration_output_1_25, A1=>nx6482, B0=>nx6462, B1=>
      nx18307);
   ix6473 : nor02_2x port map ( Y=>nx6472, A0=>data_in(25), A1=>nx35374);
   ix35401 : xnor2 port map ( Y=>nx35400, A0=>nx6510, A1=>nx18311);
   ix6511 : oai22 port map ( Y=>nx6510, A0=>nx35388, A1=>nx35403, B0=>
      nx35414, B1=>nx42571);
   ix35406 : aoi32 port map ( Y=>nx35405, A0=>nx6492, A1=>nx41931, A2=>
      nx35410, B0=>data_in(26), B1=>nx41927);
   ix6493 : nand02 port map ( Y=>nx6492, A0=>nx35408, A1=>data_in(26));
   ix35411 : nand02 port map ( Y=>nx35410, A0=>nx35412, A1=>nx6472);
   ix35413 : inv01 port map ( Y=>nx35412, A=>data_in(26));
   booth_booth_integrtaion_1_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_26, QB=>nx35414, D=>nx23281, CLK=>clk, 
      R=>rst);
   ix23272 : oai21 port map ( Y=>nx23271, A0=>nx35419, A1=>nx42553, B0=>
      nx35421);
   booth_booth_integrtaion_1_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_27, QB=>nx35419, D=>nx23271, CLK=>clk, 
      R=>rst);
   ix35422 : nand03 port map ( Y=>nx35421, A0=>nx43229, A1=>nx6654, A2=>
      nx42555);
   ix6655 : xnor2 port map ( Y=>nx6654, A0=>nx35424, A1=>nx18313);
   ix35425 : aoi22 port map ( Y=>nx35424, A0=>
      booth_booth_integration_output_1_27, A1=>nx6530, B0=>nx6510, B1=>
      nx18311);
   ix6521 : nor02_2x port map ( Y=>nx6520, A0=>data_in(27), A1=>nx35410);
   ix35437 : xnor2 port map ( Y=>nx35436, A0=>nx6558, A1=>nx18315);
   ix6559 : oai22 port map ( Y=>nx6558, A0=>nx35424, A1=>nx35439, B0=>
      nx35450, B1=>nx42573);
   ix35442 : aoi32 port map ( Y=>nx35441, A0=>nx6540, A1=>nx41933, A2=>
      nx35446, B0=>data_in(28), B1=>nx41927);
   ix6541 : nand02 port map ( Y=>nx6540, A0=>nx35444, A1=>data_in(28));
   ix35447 : nand02 port map ( Y=>nx35446, A0=>nx35448, A1=>nx6520);
   ix35449 : inv01 port map ( Y=>nx35448, A=>data_in(28));
   booth_booth_integrtaion_1_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12118, QB=>nx35450, D=>nx23261, CLK=>clk, R=>rst);
   ix23252 : oai21 port map ( Y=>nx23251, A0=>nx35455, A1=>nx42553, B0=>
      nx35457);
   booth_booth_integrtaion_1_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12117, QB=>nx35455, D=>nx23251, CLK=>clk, R=>rst);
   ix35458 : nand03 port map ( Y=>nx35457, A0=>nx43229, A1=>nx6630, A2=>
      nx42553);
   ix6631 : xnor2 port map ( Y=>nx6630, A0=>nx35460, A1=>nx18317);
   ix35461 : aoi22 port map ( Y=>nx35460, A0=>booth_output_29_dup_12117, A1
      =>nx6578, B0=>nx6558, B1=>nx18315);
   ix6569 : nor02_2x port map ( Y=>nx6568, A0=>data_in(29), A1=>nx35446);
   ix23242 : oai21 port map ( Y=>nx23241, A0=>nx35471, A1=>nx42553, B0=>
      nx35473);
   booth_booth_integrtaion_1_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx35471, D=>nx23241, CLK=>clk, R=>rst);
   ix35474 : nand03 port map ( Y=>nx35473, A0=>nx43229, A1=>nx6618, A2=>
      nx42553);
   ix6619 : xnor2 port map ( Y=>nx6618, A0=>nx6606, A1=>nx35488);
   ix6607 : oai22 port map ( Y=>nx6606, A0=>nx35460, A1=>nx35477, B0=>
      nx35471, B1=>nx42575);
   ix35480 : aoi32 port map ( Y=>nx35479, A0=>nx6588, A1=>nx41933, A2=>
      nx35484, B0=>data_in(30), B1=>nx41929);
   ix6589 : nand02 port map ( Y=>nx6588, A0=>nx35482, A1=>data_in(30));
   ix35485 : nand02 port map ( Y=>nx35484, A0=>nx35486, A1=>nx6568);
   ix35487 : inv01 port map ( Y=>nx35486, A=>data_in(30));
   ix6615 : oai22 port map ( Y=>nx6614, A0=>nx35244, A1=>nx35491, B0=>
      nx35493, B1=>nx35249);
   ix35492 : xnor2 port map ( Y=>nx35491, A0=>data_in(31), A1=>nx35484);
   ix35494 : inv01 port map ( Y=>nx35493, A=>data_in(31));
   ix35496 : aoi32 port map ( Y=>nx35495, A0=>nx6564, A1=>nx41933, A2=>
      nx35482, B0=>data_in(29), B1=>nx41929);
   ix6565 : nand02 port map ( Y=>nx6564, A0=>nx35446, A1=>data_in(29));
   ix35499 : aoi32 port map ( Y=>nx35498, A0=>nx6516, A1=>nx41933, A2=>
      nx35444, B0=>data_in(27), B1=>nx41929);
   ix6517 : nand02 port map ( Y=>nx6516, A0=>nx35410, A1=>data_in(27));
   ix35502 : aoi32 port map ( Y=>nx35501, A0=>nx6468, A1=>nx41933, A2=>
      nx35408, B0=>data_in(25), B1=>nx41929);
   ix6469 : nand02 port map ( Y=>nx6468, A0=>nx35374, A1=>data_in(25));
   ix35505 : aoi32 port map ( Y=>nx35504, A0=>nx6420, A1=>nx41933, A2=>
      nx35372, B0=>data_in(23), B1=>nx41929);
   ix6421 : nand02 port map ( Y=>nx6420, A0=>nx35338, A1=>data_in(23));
   ix35508 : aoi32 port map ( Y=>nx35507, A0=>nx6372, A1=>nx41935, A2=>
      nx35336, B0=>data_in(21), B1=>nx41929);
   ix6373 : nand02 port map ( Y=>nx6372, A0=>nx35302, A1=>data_in(21));
   ix35511 : aoi32 port map ( Y=>nx35510, A0=>nx6274, A1=>nx41935, A2=>
      nx35513, B0=>data_in(17), B1=>nx41929);
   ix6275 : nand02 port map ( Y=>nx6274, A0=>data_in(17), A1=>data_in(16));
   booth_booth_integrtaion_1_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_16, QB=>nx35224, D=>nx23381, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_15, QB=>nx35517, D=>nx23391, CLK=>clk, 
      R=>rst);
   ix6855 : aoi21 port map ( Y=>nx6854, A0=>label_2_output_0, A1=>
      booth_booth_integration_output_1_12, B0=>nx43519);
   labelsregfile_label2_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_2_output_1, QB=>nx35534, D=>nx23461, CLK=>clk, R=>rst);
   lat_label_2_input_1 : latch port map ( Q=>label_2_input_1, D=>nx6892, CLK
      =>nx41675);
   reg_label_2_input_state_machine_1 : dffr port map ( Q=>
      label_2_input_state_machine_1, QB=>OPEN, D=>nx23451, CLK=>clk, R=>rst
   );
   ix6889 : xor2 port map ( Y=>nx6888, A0=>nx35075, A1=>nx35524);
   ix35536 : xnor2 port map ( Y=>nx35535, A0=>
      booth_booth_integration_output_1_14, A1=>label_2_output_2);
   labelsregfile_label2_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_2_output_3, QB=>nx35549, D=>nx23501, CLK=>clk, R=>rst);
   lat_label_2_input_3 : latch port map ( Q=>label_2_input_3, D=>nx6956, CLK
      =>nx41675);
   reg_label_2_input_state_machine_3 : dffr port map ( Q=>
      label_2_input_state_machine_3, QB=>OPEN, D=>nx23491, CLK=>clk, R=>rst
   );
   ix6953 : xor2 port map ( Y=>nx6952, A0=>nx35064, A1=>nx35539);
   labelsregfile_label2_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_2_output_5, QB=>nx35564, D=>nx23541, CLK=>clk, R=>rst);
   lat_label_2_input_5 : latch port map ( Q=>label_2_input_5, D=>nx7020, CLK
      =>nx41675);
   reg_label_2_input_state_machine_5 : dffr port map ( Q=>
      label_2_input_state_machine_5, QB=>OPEN, D=>nx23531, CLK=>clk, R=>rst
   );
   ix7017 : xor2 port map ( Y=>nx7016, A0=>nx35053, A1=>nx35554);
   labelsregfile_label2_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_2_output_7, QB=>nx35579, D=>nx23581, CLK=>clk, R=>rst);
   lat_label_2_input_7 : latch port map ( Q=>label_2_input_7, D=>nx7084, CLK
      =>nx41675);
   reg_label_2_input_state_machine_7 : dffr port map ( Q=>
      label_2_input_state_machine_7, QB=>OPEN, D=>nx23571, CLK=>clk, R=>rst
   );
   ix7081 : xor2 port map ( Y=>nx7080, A0=>nx35042, A1=>nx35569);
   labelsregfile_label2_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_2_output_9, QB=>nx35594, D=>nx23621, CLK=>clk, R=>rst);
   lat_label_2_input_9 : latch port map ( Q=>label_2_input_9, D=>nx7148, CLK
      =>nx41677);
   reg_label_2_input_state_machine_9 : dffr port map ( Q=>
      label_2_input_state_machine_9, QB=>OPEN, D=>nx23611, CLK=>clk, R=>rst
   );
   ix7145 : xor2 port map ( Y=>nx7144, A0=>nx35031, A1=>nx35584);
   labelsregfile_label2_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_2_output_11, QB=>nx35609, D=>nx23661, CLK=>clk, R=>rst);
   lat_label_2_input_11 : latch port map ( Q=>label_2_input_11, D=>nx7212, 
      CLK=>nx41677);
   reg_label_2_input_state_machine_11 : dffr port map ( Q=>
      label_2_input_state_machine_11, QB=>OPEN, D=>nx23651, CLK=>clk, R=>rst
   );
   ix7209 : xor2 port map ( Y=>nx7208, A0=>nx35020, A1=>nx35599);
   labelsregfile_label2_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_2_output_13, QB=>nx35624, D=>nx23701, CLK=>clk, R=>rst);
   lat_label_2_input_13 : latch port map ( Q=>label_2_input_13, D=>nx7276, 
      CLK=>nx41677);
   reg_label_2_input_state_machine_13 : dffr port map ( Q=>
      label_2_input_state_machine_13, QB=>OPEN, D=>nx23691, CLK=>clk, R=>rst
   );
   ix7273 : xor2 port map ( Y=>nx7272, A0=>nx35009, A1=>nx35614);
   max_calc_reg_ans2_14 : dff port map ( Q=>max_calc_ans2_14, QB=>OPEN, D=>
      nx30101, CLK=>clk);
   ix26582 : oai21 port map ( Y=>nx26581, A0=>nx35633, A1=>nx41605, B0=>
      nx35635);
   max_calc_reg_comparator_second_inp1_14 : dff port map ( Q=>
      max_calc_comparator_second_inp1_14, QB=>nx35633, D=>nx26581, CLK=>clk
   );
   ix35636 : nand03 port map ( Y=>nx35635, A0=>nx42819, A1=>nx11808, A2=>
      nx41623);
   labelsregfile_label3_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_3_output_14, QB=>OPEN, D=>nx24541, CLK=>clk, R=>rst);
   lat_label_3_input_14 : latch port map ( Q=>label_3_input_14, D=>nx8612, 
      CLK=>nx41683);
   reg_label_3_input_state_machine_14 : dffr port map ( Q=>
      label_3_input_state_machine_14, QB=>OPEN, D=>nx23721, CLK=>clk, R=>rst
   );
   ix8609 : xnor2 port map ( Y=>nx8608, A0=>nx8604, A1=>nx36263);
   ix8605 : oai22 port map ( Y=>nx8604, A0=>nx35647, A1=>nx36252, B0=>
      nx36262, B1=>nx36021);
   ix35648 : aoi22 port map ( Y=>nx35647, A0=>label_3_output_12, A1=>
      booth_booth_integration_output_2_24, B0=>nx8540, B1=>nx18376);
   labelsregfile_label3_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_3_output_12, QB=>OPEN, D=>nx24511, CLK=>clk, R=>rst);
   lat_label_3_input_12 : latch port map ( Q=>label_3_input_12, D=>nx8554, 
      CLK=>nx41681);
   reg_label_3_input_state_machine_12 : dffr port map ( Q=>
      label_3_input_state_machine_12, QB=>OPEN, D=>nx24501, CLK=>clk, R=>rst
   );
   ix8551 : xnor2 port map ( Y=>nx8550, A0=>nx8540, A1=>nx36248);
   ix8541 : oai22 port map ( Y=>nx8540, A0=>nx35658, A1=>nx36237, B0=>
      nx36247, B1=>nx35985);
   ix35659 : aoi22 port map ( Y=>nx35658, A0=>label_3_output_10, A1=>
      booth_booth_integration_output_2_22, B0=>nx8476, B1=>nx18373);
   labelsregfile_label3_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_3_output_10, QB=>OPEN, D=>nx24471, CLK=>clk, R=>rst);
   lat_label_3_input_10 : latch port map ( Q=>label_3_input_10, D=>nx8490, 
      CLK=>nx41681);
   reg_label_3_input_state_machine_10 : dffr port map ( Q=>
      label_3_input_state_machine_10, QB=>OPEN, D=>nx24461, CLK=>clk, R=>rst
   );
   ix8487 : xnor2 port map ( Y=>nx8486, A0=>nx8476, A1=>nx36233);
   ix8477 : oai22 port map ( Y=>nx8476, A0=>nx35669, A1=>nx36222, B0=>
      nx36232, B1=>nx35949);
   ix35670 : aoi22 port map ( Y=>nx35669, A0=>label_3_output_8, A1=>
      booth_booth_integration_output_2_20, B0=>nx8412, B1=>nx18369);
   labelsregfile_label3_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_3_output_8, QB=>OPEN, D=>nx24431, CLK=>clk, R=>rst);
   lat_label_3_input_8 : latch port map ( Q=>label_3_input_8, D=>nx8426, CLK
      =>nx41681);
   reg_label_3_input_state_machine_8 : dffr port map ( Q=>
      label_3_input_state_machine_8, QB=>OPEN, D=>nx24421, CLK=>clk, R=>rst
   );
   ix8423 : xnor2 port map ( Y=>nx8422, A0=>nx8412, A1=>nx36218);
   ix8413 : oai22 port map ( Y=>nx8412, A0=>nx35680, A1=>nx36207, B0=>
      nx36217, B1=>nx35911);
   ix35681 : aoi22 port map ( Y=>nx35680, A0=>label_3_output_6, A1=>
      booth_booth_integration_output_2_18, B0=>nx8348, B1=>nx18367);
   labelsregfile_label3_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_3_output_6, QB=>OPEN, D=>nx24391, CLK=>clk, R=>rst);
   lat_label_3_input_6 : latch port map ( Q=>label_3_input_6, D=>nx8362, CLK
      =>nx41679);
   reg_label_3_input_state_machine_6 : dffr port map ( Q=>
      label_3_input_state_machine_6, QB=>OPEN, D=>nx24381, CLK=>clk, R=>rst
   );
   ix8359 : xnor2 port map ( Y=>nx8358, A0=>nx8348, A1=>nx36203);
   ix8349 : oai22 port map ( Y=>nx8348, A0=>nx35691, A1=>nx36192, B0=>
      nx36202, B1=>nx35872);
   ix35692 : aoi22 port map ( Y=>nx35691, A0=>label_3_output_4, A1=>
      booth_booth_integration_output_2_16, B0=>nx8284, B1=>nx18365);
   labelsregfile_label3_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_3_output_4, QB=>OPEN, D=>nx24351, CLK=>clk, R=>rst);
   lat_label_3_input_4 : latch port map ( Q=>label_3_input_4, D=>nx8298, CLK
      =>nx41679);
   reg_label_3_input_state_machine_4 : dffr port map ( Q=>
      label_3_input_state_machine_4, QB=>OPEN, D=>nx24341, CLK=>clk, R=>rst
   );
   ix8295 : xnor2 port map ( Y=>nx8294, A0=>nx8284, A1=>nx36188);
   ix8285 : oai22 port map ( Y=>nx8284, A0=>nx35702, A1=>nx36177, B0=>
      nx36187, B1=>nx36155);
   ix35703 : aoi22 port map ( Y=>nx35702, A0=>label_3_output_2, A1=>
      booth_booth_integration_output_2_14, B0=>nx8220, B1=>nx18363);
   labelsregfile_label3_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_3_output_2, QB=>OPEN, D=>nx24311, CLK=>clk, R=>rst);
   lat_label_3_input_2 : latch port map ( Q=>label_3_input_2, D=>nx8234, CLK
      =>nx41679);
   reg_label_3_input_state_machine_2 : dffr port map ( Q=>
      label_3_input_state_machine_2, QB=>OPEN, D=>nx24301, CLK=>clk, R=>rst
   );
   ix8231 : xnor2 port map ( Y=>nx8230, A0=>nx8220, A1=>nx36173);
   ix8221 : oai22 port map ( Y=>nx8220, A0=>nx35713, A1=>nx36162, B0=>
      nx36172, B1=>nx36158);
   ix35714 : nand02 port map ( Y=>nx35713, A0=>label_3_output_0, A1=>
      booth_booth_integration_output_2_12);
   labelsregfile_label3_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_3_output_0, QB=>OPEN, D=>nx24271, CLK=>clk, R=>rst);
   lat_label_3_input_0 : latch port map ( Q=>label_3_input_0, D=>nx8176, CLK
      =>nx41679);
   ix8177 : oai21 port map ( Y=>nx8176, A0=>nx35719, A1=>nx41439, B0=>
      nx35723);
   reg_label_3_input_state_machine_0 : dffr port map ( Q=>
      label_3_input_state_machine_0, QB=>nx35719, D=>nx24261, CLK=>clk, R=>
      rst);
   ix35724 : oai21 port map ( Y=>nx35723, A0=>
      booth_booth_integration_output_2_12, A1=>label_3_output_0, B0=>nx8164
   );
   booth_booth_integrtaion_2_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_12, QB=>OPEN, D=>nx24251, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_13, QB=>nx36158, D=>nx24241, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_14, QB=>OPEN, D=>nx24231, CLK=>clk, R
      =>rst);
   ix35737 : aoi22 port map ( Y=>nx35736, A0=>nx41795, A1=>nx41951, B0=>
      nx8106, B1=>nx8112);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_reg_output_0, QB=>OPEN, 
      D=>nx23751, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_0, QB=>OPEN, D=>nx23737, CLK
      =>clk, S=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_reg_output_9, QB=>OPEN, 
      D=>nx23931, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_9, QB=>OPEN, D=>nx23921, CLK
      =>clk, R=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12744, QB=>OPEN, D=>nx23911, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_8, QB=>OPEN, D=>nx23901, CLK
      =>clk, R=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12745, QB=>OPEN, D=>nx23891, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_7, QB=>OPEN, D=>nx23881, CLK
      =>clk, R=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12746, QB=>OPEN, D=>nx23871, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_6, QB=>OPEN, D=>nx23861, CLK
      =>clk, R=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12747, QB=>OPEN, D=>nx23851, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_5, QB=>OPEN, D=>nx23841, CLK
      =>clk, R=>nx41489);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12748, QB=>OPEN, D=>nx23831, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_4, QB=>OPEN, D=>nx23821, CLK
      =>clk, R=>nx41487);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12749, QB=>OPEN, D=>nx23811, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_3, QB=>OPEN, D=>nx23801, CLK
      =>clk, R=>nx41487);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12750, QB=>OPEN, D=>nx23791, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_2, QB=>OPEN, D=>nx23781, CLK
      =>clk, R=>nx41487);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12751, QB=>OPEN, D=>nx23771, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_1, QB=>OPEN, D=>nx23761, CLK
      =>clk, R=>nx41487);
   ix23732 : nand02 port map ( Y=>nx23731, A0=>nx42941, A1=>nx41937);
   booth_booth_integrtaion_2_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx35783, D=>nx23731, CLK=>clk, S=>nx41487);
   ix8107 : nand02 port map ( Y=>nx8106, A0=>nx35804, A1=>nx35862);
   ix35805 : oai21 port map ( Y=>nx35804, A0=>nx41963, A1=>nx41959, B0=>
      data_in(32));
   ix24062 : oai21 port map ( Y=>nx24061, A0=>nx35809, A1=>nx42577, B0=>
      nx35811);
   booth_booth_integrtaion_2_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx35809, D=>nx24061, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12149, QB=>nx35860, D=>nx24051, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12148, QB=>OPEN, D=>nx24041, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12147, QB=>OPEN, D=>nx24031, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12146, QB=>OPEN, D=>nx24021, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12145, QB=>OPEN, D=>nx24011, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12144, QB=>OPEN, D=>nx24001, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12143, QB=>OPEN, D=>nx23991, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12142, QB=>OPEN, D=>nx23981, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12141, QB=>OPEN, D=>nx23971, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12140, QB=>OPEN, D=>nx23961, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12139, QB=>OPEN, D=>nx23951, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12138, QB=>OPEN, D=>nx23941, CLK=>clk, R=>rst);
   ix35867 : xnor2 port map ( Y=>nx35866, A0=>nx7576, A1=>nx18337);
   ix24202 : oai21 port map ( Y=>nx24201, A0=>nx35872, A1=>nx42577, B0=>
      nx35874);
   booth_booth_integrtaion_2_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_17, QB=>nx35872, D=>nx24201, CLK=>clk, 
      R=>rst);
   ix35875 : nand03 port map ( Y=>nx35874, A0=>nx42585, A1=>nx8084, A2=>
      nx42581);
   ix8085 : xnor2 port map ( Y=>nx8084, A0=>nx35877, A1=>nx18339);
   ix35878 : aoi22 port map ( Y=>nx35877, A0=>
      booth_booth_integration_output_2_17, A1=>nx7600, B0=>nx7576, B1=>
      nx18337);
   ix7591 : nor02_2x port map ( Y=>nx7590, A0=>data_in(32), A1=>data_in(33)
   );
   ix24192 : oai21 port map ( Y=>nx24191, A0=>nx35892, A1=>nx42577, B0=>
      nx35894);
   booth_booth_integrtaion_2_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_18, QB=>nx35892, D=>nx24191, CLK=>clk, 
      R=>rst);
   ix35895 : nand03 port map ( Y=>nx35894, A0=>nx42585, A1=>nx8072, A2=>
      nx42581);
   ix8073 : xnor2 port map ( Y=>nx8072, A0=>nx7628, A1=>nx35907);
   ix7629 : oai22 port map ( Y=>nx7628, A0=>nx35877, A1=>nx35898, B0=>
      nx35892, B1=>nx42589);
   ix35901 : aoi32 port map ( Y=>nx35900, A0=>nx7610, A1=>nx41963, A2=>
      nx35903, B0=>data_in(34), B1=>nx41959);
   ix7611 : oai21 port map ( Y=>nx7610, A0=>data_in(32), A1=>data_in(33), B0
      =>data_in(34));
   ix24182 : oai21 port map ( Y=>nx24181, A0=>nx35911, A1=>nx42577, B0=>
      nx35913);
   booth_booth_integrtaion_2_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_19, QB=>nx35911, D=>nx24181, CLK=>clk, 
      R=>rst);
   ix35914 : nand03 port map ( Y=>nx35913, A0=>nx42585, A1=>nx8060, A2=>
      nx42581);
   ix8061 : xnor2 port map ( Y=>nx8060, A0=>nx35916, A1=>nx18343);
   ix35917 : aoi22 port map ( Y=>nx35916, A0=>
      booth_booth_integration_output_2_19, A1=>nx7648, B0=>nx7628, B1=>
      nx18341);
   ix7649 : oai32 port map ( Y=>nx7648, A0=>nx35919, A1=>nx35882, A2=>nx7638, 
      B0=>nx35922, B1=>nx35887);
   ix7615 : nor03_2x port map ( Y=>nx7614, A0=>data_in(34), A1=>data_in(32), 
      A2=>data_in(33));
   ix35923 : inv01 port map ( Y=>nx35922, A=>data_in(35));
   ix7639 : nor04 port map ( Y=>nx7638, A0=>data_in(35), A1=>data_in(34), A2
      =>data_in(32), A3=>data_in(33));
   ix35931 : xnor2 port map ( Y=>nx35930, A0=>nx7676, A1=>nx18345);
   ix7677 : oai22 port map ( Y=>nx7676, A0=>nx35916, A1=>nx35933, B0=>
      nx35944, B1=>nx42591);
   ix35936 : aoi32 port map ( Y=>nx35935, A0=>nx7658, A1=>nx41963, A2=>
      nx35940, B0=>data_in(36), B1=>nx41959);
   ix7659 : nand02 port map ( Y=>nx7658, A0=>nx35938, A1=>data_in(36));
   ix35941 : nand02 port map ( Y=>nx35940, A0=>nx35942, A1=>nx7638);
   ix35943 : inv01 port map ( Y=>nx35942, A=>data_in(36));
   booth_booth_integrtaion_2_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_20, QB=>nx35944, D=>nx24171, CLK=>clk, 
      R=>rst);
   ix24162 : oai21 port map ( Y=>nx24161, A0=>nx35949, A1=>nx42577, B0=>
      nx35951);
   booth_booth_integrtaion_2_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_21, QB=>nx35949, D=>nx24161, CLK=>clk, 
      R=>rst);
   ix35952 : nand03 port map ( Y=>nx35951, A0=>nx42585, A1=>nx8036, A2=>
      nx42581);
   ix8037 : xnor2 port map ( Y=>nx8036, A0=>nx35954, A1=>nx18347);
   ix35955 : aoi22 port map ( Y=>nx35954, A0=>
      booth_booth_integration_output_2_21, A1=>nx7696, B0=>nx7676, B1=>
      nx18345);
   ix7687 : nor02_2x port map ( Y=>nx7686, A0=>data_in(37), A1=>nx35940);
   ix35967 : xnor2 port map ( Y=>nx35966, A0=>nx7724, A1=>nx18349);
   ix7725 : oai22 port map ( Y=>nx7724, A0=>nx35954, A1=>nx35969, B0=>
      nx35980, B1=>nx42593);
   ix35972 : aoi32 port map ( Y=>nx35971, A0=>nx7706, A1=>nx41963, A2=>
      nx35976, B0=>data_in(38), B1=>nx41959);
   ix7707 : nand02 port map ( Y=>nx7706, A0=>nx35974, A1=>data_in(38));
   ix35977 : nand02 port map ( Y=>nx35976, A0=>nx35978, A1=>nx7686);
   ix35979 : inv01 port map ( Y=>nx35978, A=>data_in(38));
   booth_booth_integrtaion_2_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_22, QB=>nx35980, D=>nx24151, CLK=>clk, 
      R=>rst);
   ix24142 : oai21 port map ( Y=>nx24141, A0=>nx35985, A1=>nx42579, B0=>
      nx35987);
   booth_booth_integrtaion_2_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_23, QB=>nx35985, D=>nx24141, CLK=>clk, 
      R=>rst);
   ix35988 : nand03 port map ( Y=>nx35987, A0=>nx42585, A1=>nx8012, A2=>
      nx42581);
   ix8013 : xnor2 port map ( Y=>nx8012, A0=>nx35990, A1=>nx18350);
   ix35991 : aoi22 port map ( Y=>nx35990, A0=>
      booth_booth_integration_output_2_23, A1=>nx7744, B0=>nx7724, B1=>
      nx18349);
   ix7735 : nor02_2x port map ( Y=>nx7734, A0=>data_in(39), A1=>nx35976);
   ix36003 : xnor2 port map ( Y=>nx36002, A0=>nx7772, A1=>nx18351);
   ix7773 : oai22 port map ( Y=>nx7772, A0=>nx35990, A1=>nx36005, B0=>
      nx36016, B1=>nx42595);
   ix36008 : aoi32 port map ( Y=>nx36007, A0=>nx7754, A1=>nx41963, A2=>
      nx36012, B0=>data_in(40), B1=>nx41959);
   ix7755 : nand02 port map ( Y=>nx7754, A0=>nx36010, A1=>data_in(40));
   ix36013 : nand02 port map ( Y=>nx36012, A0=>nx36014, A1=>nx7734);
   ix36015 : inv01 port map ( Y=>nx36014, A=>data_in(40));
   booth_booth_integrtaion_2_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_24, QB=>nx36016, D=>nx24131, CLK=>clk, 
      R=>rst);
   ix24122 : oai21 port map ( Y=>nx24121, A0=>nx36021, A1=>nx42579, B0=>
      nx36023);
   booth_booth_integrtaion_2_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_25, QB=>nx36021, D=>nx24121, CLK=>clk, 
      R=>rst);
   ix36024 : nand03 port map ( Y=>nx36023, A0=>nx42585, A1=>nx7988, A2=>
      nx42581);
   ix7989 : xnor2 port map ( Y=>nx7988, A0=>nx36026, A1=>nx18352);
   ix36027 : aoi22 port map ( Y=>nx36026, A0=>
      booth_booth_integration_output_2_25, A1=>nx7792, B0=>nx7772, B1=>
      nx18351);
   ix7783 : nor02_2x port map ( Y=>nx7782, A0=>data_in(41), A1=>nx36012);
   ix36039 : xnor2 port map ( Y=>nx36038, A0=>nx7820, A1=>nx18353);
   ix7821 : oai22 port map ( Y=>nx7820, A0=>nx36026, A1=>nx36041, B0=>
      nx36052, B1=>nx42597);
   ix36044 : aoi32 port map ( Y=>nx36043, A0=>nx7802, A1=>nx41963, A2=>
      nx36048, B0=>data_in(42), B1=>nx41959);
   ix7803 : nand02 port map ( Y=>nx7802, A0=>nx36046, A1=>data_in(42));
   ix36049 : nand02 port map ( Y=>nx36048, A0=>nx36050, A1=>nx7782);
   ix36051 : inv01 port map ( Y=>nx36050, A=>data_in(42));
   booth_booth_integrtaion_2_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_26, QB=>nx36052, D=>nx24111, CLK=>clk, 
      R=>rst);
   ix24102 : oai21 port map ( Y=>nx24101, A0=>nx36057, A1=>nx42579, B0=>
      nx36059);
   booth_booth_integrtaion_2_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_27, QB=>nx36057, D=>nx24101, CLK=>clk, 
      R=>rst);
   ix36060 : nand03 port map ( Y=>nx36059, A0=>nx43243, A1=>nx7964, A2=>
      nx42581);
   ix7965 : xnor2 port map ( Y=>nx7964, A0=>nx36062, A1=>nx18354);
   ix36063 : aoi22 port map ( Y=>nx36062, A0=>
      booth_booth_integration_output_2_27, A1=>nx7840, B0=>nx7820, B1=>
      nx18353);
   ix7831 : nor02_2x port map ( Y=>nx7830, A0=>data_in(43), A1=>nx36048);
   ix36075 : xnor2 port map ( Y=>nx36074, A0=>nx7868, A1=>nx18355);
   ix7869 : oai22 port map ( Y=>nx7868, A0=>nx36062, A1=>nx36077, B0=>
      nx36088, B1=>nx42599);
   ix36080 : aoi32 port map ( Y=>nx36079, A0=>nx7850, A1=>nx41965, A2=>
      nx36084, B0=>data_in(44), B1=>nx41959);
   ix7851 : nand02 port map ( Y=>nx7850, A0=>nx36082, A1=>data_in(44));
   ix36085 : nand02 port map ( Y=>nx36084, A0=>nx36086, A1=>nx7830);
   ix36087 : inv01 port map ( Y=>nx36086, A=>data_in(44));
   booth_booth_integrtaion_2_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12137, QB=>nx36088, D=>nx24091, CLK=>clk, R=>rst);
   ix24082 : oai21 port map ( Y=>nx24081, A0=>nx36093, A1=>nx42579, B0=>
      nx36095);
   booth_booth_integrtaion_2_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12136, QB=>nx36093, D=>nx24081, CLK=>clk, R=>rst);
   ix36096 : nand03 port map ( Y=>nx36095, A0=>nx43243, A1=>nx7940, A2=>
      nx42579);
   ix7941 : xnor2 port map ( Y=>nx7940, A0=>nx36098, A1=>nx18357);
   ix36099 : aoi22 port map ( Y=>nx36098, A0=>booth_output_29_dup_12136, A1
      =>nx7888, B0=>nx7868, B1=>nx18355);
   ix7879 : nor02_2x port map ( Y=>nx7878, A0=>data_in(45), A1=>nx36084);
   ix24072 : oai21 port map ( Y=>nx24071, A0=>nx36109, A1=>nx42579, B0=>
      nx36111);
   booth_booth_integrtaion_2_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx36109, D=>nx24071, CLK=>clk, R=>rst);
   ix36112 : nand03 port map ( Y=>nx36111, A0=>nx43243, A1=>nx7928, A2=>
      nx42579);
   ix7929 : xnor2 port map ( Y=>nx7928, A0=>nx7916, A1=>nx36126);
   ix7917 : oai22 port map ( Y=>nx7916, A0=>nx36098, A1=>nx36115, B0=>
      nx36109, B1=>nx42601);
   ix36118 : aoi32 port map ( Y=>nx36117, A0=>nx7898, A1=>nx41965, A2=>
      nx36122, B0=>data_in(46), B1=>nx41961);
   ix7899 : nand02 port map ( Y=>nx7898, A0=>nx36120, A1=>data_in(46));
   ix36123 : nand02 port map ( Y=>nx36122, A0=>nx36124, A1=>nx7878);
   ix36125 : inv01 port map ( Y=>nx36124, A=>data_in(46));
   ix7925 : oai22 port map ( Y=>nx7924, A0=>nx35882, A1=>nx36129, B0=>
      nx36131, B1=>nx35887);
   ix36130 : xnor2 port map ( Y=>nx36129, A0=>data_in(47), A1=>nx36122);
   ix36132 : inv01 port map ( Y=>nx36131, A=>data_in(47));
   ix36134 : aoi32 port map ( Y=>nx36133, A0=>nx7874, A1=>nx41965, A2=>
      nx36120, B0=>data_in(45), B1=>nx41961);
   ix7875 : nand02 port map ( Y=>nx7874, A0=>nx36084, A1=>data_in(45));
   ix36137 : aoi32 port map ( Y=>nx36136, A0=>nx7826, A1=>nx41965, A2=>
      nx36082, B0=>data_in(43), B1=>nx41961);
   ix7827 : nand02 port map ( Y=>nx7826, A0=>nx36048, A1=>data_in(43));
   ix36140 : aoi32 port map ( Y=>nx36139, A0=>nx7778, A1=>nx41965, A2=>
      nx36046, B0=>data_in(41), B1=>nx41961);
   ix7779 : nand02 port map ( Y=>nx7778, A0=>nx36012, A1=>data_in(41));
   ix36143 : aoi32 port map ( Y=>nx36142, A0=>nx7730, A1=>nx41965, A2=>
      nx36010, B0=>data_in(39), B1=>nx41961);
   ix7731 : nand02 port map ( Y=>nx7730, A0=>nx35976, A1=>data_in(39));
   ix36146 : aoi32 port map ( Y=>nx36145, A0=>nx7682, A1=>nx41967, A2=>
      nx35974, B0=>data_in(37), B1=>nx41961);
   ix7683 : nand02 port map ( Y=>nx7682, A0=>nx35940, A1=>data_in(37));
   ix36149 : aoi32 port map ( Y=>nx36148, A0=>nx7584, A1=>nx41967, A2=>
      nx36151, B0=>data_in(33), B1=>nx41961);
   ix7585 : nand02 port map ( Y=>nx7584, A0=>data_in(33), A1=>data_in(32));
   booth_booth_integrtaion_2_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_16, QB=>nx35862, D=>nx24211, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_15, QB=>nx36155, D=>nx24221, CLK=>clk, 
      R=>rst);
   ix8165 : aoi21 port map ( Y=>nx8164, A0=>label_3_output_0, A1=>
      booth_booth_integration_output_2_12, B0=>nx43519);
   labelsregfile_label3_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_3_output_1, QB=>nx36172, D=>nx24291, CLK=>clk, R=>rst);
   lat_label_3_input_1 : latch port map ( Q=>label_3_input_1, D=>nx8202, CLK
      =>nx41679);
   reg_label_3_input_state_machine_1 : dffr port map ( Q=>
      label_3_input_state_machine_1, QB=>OPEN, D=>nx24281, CLK=>clk, R=>rst
   );
   ix8199 : xor2 port map ( Y=>nx8198, A0=>nx35713, A1=>nx36162);
   ix36174 : xnor2 port map ( Y=>nx36173, A0=>
      booth_booth_integration_output_2_14, A1=>label_3_output_2);
   labelsregfile_label3_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_3_output_3, QB=>nx36187, D=>nx24331, CLK=>clk, R=>rst);
   lat_label_3_input_3 : latch port map ( Q=>label_3_input_3, D=>nx8266, CLK
      =>nx41679);
   reg_label_3_input_state_machine_3 : dffr port map ( Q=>
      label_3_input_state_machine_3, QB=>OPEN, D=>nx24321, CLK=>clk, R=>rst
   );
   ix8263 : xor2 port map ( Y=>nx8262, A0=>nx35702, A1=>nx36177);
   labelsregfile_label3_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_3_output_5, QB=>nx36202, D=>nx24371, CLK=>clk, R=>rst);
   lat_label_3_input_5 : latch port map ( Q=>label_3_input_5, D=>nx8330, CLK
      =>nx41679);
   reg_label_3_input_state_machine_5 : dffr port map ( Q=>
      label_3_input_state_machine_5, QB=>OPEN, D=>nx24361, CLK=>clk, R=>rst
   );
   ix8327 : xor2 port map ( Y=>nx8326, A0=>nx35691, A1=>nx36192);
   labelsregfile_label3_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_3_output_7, QB=>nx36217, D=>nx24411, CLK=>clk, R=>rst);
   lat_label_3_input_7 : latch port map ( Q=>label_3_input_7, D=>nx8394, CLK
      =>nx41681);
   reg_label_3_input_state_machine_7 : dffr port map ( Q=>
      label_3_input_state_machine_7, QB=>OPEN, D=>nx24401, CLK=>clk, R=>rst
   );
   ix8391 : xor2 port map ( Y=>nx8390, A0=>nx35680, A1=>nx36207);
   labelsregfile_label3_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_3_output_9, QB=>nx36232, D=>nx24451, CLK=>clk, R=>rst);
   lat_label_3_input_9 : latch port map ( Q=>label_3_input_9, D=>nx8458, CLK
      =>nx41681);
   reg_label_3_input_state_machine_9 : dffr port map ( Q=>
      label_3_input_state_machine_9, QB=>OPEN, D=>nx24441, CLK=>clk, R=>rst
   );
   ix8455 : xor2 port map ( Y=>nx8454, A0=>nx35669, A1=>nx36222);
   labelsregfile_label3_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_3_output_11, QB=>nx36247, D=>nx24491, CLK=>clk, R=>rst);
   lat_label_3_input_11 : latch port map ( Q=>label_3_input_11, D=>nx8522, 
      CLK=>nx41681);
   reg_label_3_input_state_machine_11 : dffr port map ( Q=>
      label_3_input_state_machine_11, QB=>OPEN, D=>nx24481, CLK=>clk, R=>rst
   );
   ix8519 : xor2 port map ( Y=>nx8518, A0=>nx35658, A1=>nx36237);
   labelsregfile_label3_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_3_output_13, QB=>nx36262, D=>nx24531, CLK=>clk, R=>rst);
   lat_label_3_input_13 : latch port map ( Q=>label_3_input_13, D=>nx8586, 
      CLK=>nx41681);
   reg_label_3_input_state_machine_13 : dffr port map ( Q=>
      label_3_input_state_machine_13, QB=>OPEN, D=>nx24521, CLK=>clk, R=>rst
   );
   ix8583 : xor2 port map ( Y=>nx8582, A0=>nx35647, A1=>nx36252);
   max_calc_reg_ans3_14 : dff port map ( Q=>max_calc_ans3_14, QB=>OPEN, D=>
      nx26571, CLK=>clk);
   ix26572 : ao32 port map ( Y=>nx26571, A0=>nx42819, A1=>nx11794, A2=>
      nx41811, B0=>max_calc_ans3_14, B1=>nx42679);
   ix25382 : oai21 port map ( Y=>nx25381, A0=>nx36271, A1=>nx41605, B0=>
      nx36273);
   max_calc_reg_comparator_third_inp1_14 : dff port map ( Q=>
      max_calc_comparator_third_inp1_14, QB=>nx36271, D=>nx25381, CLK=>clk);
   ix36274 : nand03 port map ( Y=>nx36273, A0=>label_5_output_14, A1=>
      nx42631, A2=>nx41605);
   labelsregfile_label5_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_5_output_14, QB=>OPEN, D=>nx25371, CLK=>clk, R=>rst);
   lat_label_5_input_14 : latch port map ( Q=>label_5_input_14, D=>nx9932, 
      CLK=>nx41687);
   reg_label_5_input_state_machine_14 : dffr port map ( Q=>
      label_5_input_state_machine_14, QB=>OPEN, D=>nx24551, CLK=>clk, R=>rst
   );
   ix9929 : xnor2 port map ( Y=>nx9928, A0=>nx9924, A1=>nx36900);
   ix9925 : oai22 port map ( Y=>nx9924, A0=>nx36284, A1=>nx36889, B0=>
      nx36899, B1=>nx36658);
   ix36285 : aoi22 port map ( Y=>nx36284, A0=>label_5_output_12, A1=>
      booth_booth_integration_output_4_24, B0=>nx9860, B1=>nx18415);
   labelsregfile_label5_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_5_output_12, QB=>OPEN, D=>nx25341, CLK=>clk, R=>rst);
   lat_label_5_input_12 : latch port map ( Q=>label_5_input_12, D=>nx9874, 
      CLK=>nx41685);
   reg_label_5_input_state_machine_12 : dffr port map ( Q=>
      label_5_input_state_machine_12, QB=>OPEN, D=>nx25331, CLK=>clk, R=>rst
   );
   ix9871 : xnor2 port map ( Y=>nx9870, A0=>nx9860, A1=>nx36885);
   ix9861 : oai22 port map ( Y=>nx9860, A0=>nx36295, A1=>nx36874, B0=>
      nx36884, B1=>nx36622);
   ix36296 : aoi22 port map ( Y=>nx36295, A0=>label_5_output_10, A1=>
      booth_booth_integration_output_4_22, B0=>nx9796, B1=>nx18411);
   labelsregfile_label5_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_5_output_10, QB=>OPEN, D=>nx25301, CLK=>clk, R=>rst);
   lat_label_5_input_10 : latch port map ( Q=>label_5_input_10, D=>nx9810, 
      CLK=>nx41685);
   reg_label_5_input_state_machine_10 : dffr port map ( Q=>
      label_5_input_state_machine_10, QB=>OPEN, D=>nx25291, CLK=>clk, R=>rst
   );
   ix9807 : xnor2 port map ( Y=>nx9806, A0=>nx9796, A1=>nx36870);
   ix9797 : oai22 port map ( Y=>nx9796, A0=>nx36306, A1=>nx36859, B0=>
      nx36869, B1=>nx36586);
   ix36307 : aoi22 port map ( Y=>nx36306, A0=>label_5_output_8, A1=>
      booth_booth_integration_output_4_20, B0=>nx9732, B1=>nx18407);
   labelsregfile_label5_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_5_output_8, QB=>OPEN, D=>nx25261, CLK=>clk, R=>rst);
   lat_label_5_input_8 : latch port map ( Q=>label_5_input_8, D=>nx9746, CLK
      =>nx41685);
   reg_label_5_input_state_machine_8 : dffr port map ( Q=>
      label_5_input_state_machine_8, QB=>OPEN, D=>nx25251, CLK=>clk, R=>rst
   );
   ix9743 : xnor2 port map ( Y=>nx9742, A0=>nx9732, A1=>nx36855);
   ix9733 : oai22 port map ( Y=>nx9732, A0=>nx36317, A1=>nx36844, B0=>
      nx36854, B1=>nx36548);
   ix36318 : aoi22 port map ( Y=>nx36317, A0=>label_5_output_6, A1=>
      booth_booth_integration_output_4_18, B0=>nx9668, B1=>nx18405);
   labelsregfile_label5_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_5_output_6, QB=>OPEN, D=>nx25221, CLK=>clk, R=>rst);
   lat_label_5_input_6 : latch port map ( Q=>label_5_input_6, D=>nx9682, CLK
      =>nx41685);
   reg_label_5_input_state_machine_6 : dffr port map ( Q=>
      label_5_input_state_machine_6, QB=>OPEN, D=>nx25211, CLK=>clk, R=>rst
   );
   ix9679 : xnor2 port map ( Y=>nx9678, A0=>nx9668, A1=>nx36840);
   ix9669 : oai22 port map ( Y=>nx9668, A0=>nx36328, A1=>nx36829, B0=>
      nx36839, B1=>nx36509);
   ix36329 : aoi22 port map ( Y=>nx36328, A0=>label_5_output_4, A1=>
      booth_booth_integration_output_4_16, B0=>nx9604, B1=>nx18403);
   labelsregfile_label5_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_5_output_4, QB=>OPEN, D=>nx25181, CLK=>clk, R=>rst);
   lat_label_5_input_4 : latch port map ( Q=>label_5_input_4, D=>nx9618, CLK
      =>nx41683);
   reg_label_5_input_state_machine_4 : dffr port map ( Q=>
      label_5_input_state_machine_4, QB=>OPEN, D=>nx25171, CLK=>clk, R=>rst
   );
   ix9615 : xnor2 port map ( Y=>nx9614, A0=>nx9604, A1=>nx36825);
   ix9605 : oai22 port map ( Y=>nx9604, A0=>nx36339, A1=>nx36814, B0=>
      nx36824, B1=>nx36792);
   ix36340 : aoi22 port map ( Y=>nx36339, A0=>label_5_output_2, A1=>
      booth_booth_integration_output_4_14, B0=>nx9540, B1=>nx18401);
   labelsregfile_label5_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_5_output_2, QB=>OPEN, D=>nx25141, CLK=>clk, R=>rst);
   lat_label_5_input_2 : latch port map ( Q=>label_5_input_2, D=>nx9554, CLK
      =>nx41683);
   reg_label_5_input_state_machine_2 : dffr port map ( Q=>
      label_5_input_state_machine_2, QB=>OPEN, D=>nx25131, CLK=>clk, R=>rst
   );
   ix9551 : xnor2 port map ( Y=>nx9550, A0=>nx9540, A1=>nx36810);
   ix9541 : oai22 port map ( Y=>nx9540, A0=>nx36350, A1=>nx36799, B0=>
      nx36809, B1=>nx36795);
   ix36351 : nand02 port map ( Y=>nx36350, A0=>label_5_output_0, A1=>
      booth_booth_integration_output_4_12);
   labelsregfile_label5_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_5_output_0, QB=>OPEN, D=>nx25101, CLK=>clk, R=>rst);
   lat_label_5_input_0 : latch port map ( Q=>label_5_input_0, D=>nx9496, CLK
      =>nx41683);
   ix9497 : oai21 port map ( Y=>nx9496, A0=>nx36356, A1=>nx41443, B0=>
      nx36360);
   reg_label_5_input_state_machine_0 : dffr port map ( Q=>
      label_5_input_state_machine_0, QB=>nx36356, D=>nx25091, CLK=>clk, R=>
      rst);
   ix36361 : oai21 port map ( Y=>nx36360, A0=>
      booth_booth_integration_output_4_12, A1=>label_5_output_0, B0=>nx9484
   );
   booth_booth_integrtaion_4_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_12, QB=>OPEN, D=>nx25081, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_13, QB=>nx36795, D=>nx25071, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_14, QB=>OPEN, D=>nx25061, CLK=>clk, R
      =>rst);
   ix36374 : aoi22 port map ( Y=>nx36373, A0=>nx41795, A1=>nx41983, B0=>
      nx9426, B1=>nx9432);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_reg_output_0, QB=>OPEN, 
      D=>nx24581, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_0, QB=>OPEN, D=>nx24567, CLK
      =>clk, S=>nx41493);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_reg_output_9, QB=>OPEN, 
      D=>nx24761, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_9, QB=>OPEN, D=>nx24751, CLK
      =>clk, R=>nx41493);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12800, QB=>OPEN, D=>nx24741, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_8, QB=>OPEN, D=>nx24731, CLK
      =>clk, R=>nx41493);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12801, QB=>OPEN, D=>nx24721, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_7, QB=>OPEN, D=>nx24711, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12802, QB=>OPEN, D=>nx24701, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_6, QB=>OPEN, D=>nx24691, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12803, QB=>OPEN, D=>nx24681, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_5, QB=>OPEN, D=>nx24671, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12804, QB=>OPEN, D=>nx24661, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_4, QB=>OPEN, D=>nx24651, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12805, QB=>OPEN, D=>nx24641, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_3, QB=>OPEN, D=>nx24631, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12806, QB=>OPEN, D=>nx24621, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_2, QB=>OPEN, D=>nx24611, CLK
      =>clk, R=>nx41491);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12807, QB=>OPEN, D=>nx24601, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_1, QB=>OPEN, D=>nx24591, CLK
      =>clk, R=>nx41489);
   ix24562 : nand02 port map ( Y=>nx24561, A0=>nx42945, A1=>nx41969);
   booth_booth_integrtaion_4_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx36420, D=>nx24561, CLK=>clk, S=>nx41491);
   ix9427 : nand02 port map ( Y=>nx9426, A0=>nx36441, A1=>nx36499);
   ix36442 : oai21 port map ( Y=>nx36441, A0=>nx41995, A1=>nx41991, B0=>
      data_in(64));
   ix24892 : oai21 port map ( Y=>nx24891, A0=>nx36446, A1=>nx42603, B0=>
      nx36448);
   booth_booth_integrtaion_4_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx36446, D=>nx24891, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12187, QB=>nx36497, D=>nx24881, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12186, QB=>OPEN, D=>nx24871, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12185, QB=>OPEN, D=>nx24861, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12184, QB=>OPEN, D=>nx24851, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12183, QB=>OPEN, D=>nx24841, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12182, QB=>OPEN, D=>nx24831, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12181, QB=>OPEN, D=>nx24821, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12180, QB=>OPEN, D=>nx24811, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12179, QB=>OPEN, D=>nx24801, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12178, QB=>OPEN, D=>nx24791, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12177, QB=>OPEN, D=>nx24781, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12176, QB=>OPEN, D=>nx24771, CLK=>clk, R=>rst);
   ix36504 : xnor2 port map ( Y=>nx36503, A0=>nx8896, A1=>nx18379);
   ix25032 : oai21 port map ( Y=>nx25031, A0=>nx36509, A1=>nx42603, B0=>
      nx36511);
   booth_booth_integrtaion_4_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_17, QB=>nx36509, D=>nx25031, CLK=>clk, 
      R=>rst);
   ix36512 : nand03 port map ( Y=>nx36511, A0=>nx42611, A1=>nx9404, A2=>
      nx42607);
   ix9405 : xnor2 port map ( Y=>nx9404, A0=>nx36514, A1=>nx18380);
   ix36515 : aoi22 port map ( Y=>nx36514, A0=>
      booth_booth_integration_output_4_17, A1=>nx8920, B0=>nx8896, B1=>
      nx18379);
   ix8911 : nor02_2x port map ( Y=>nx8910, A0=>data_in(64), A1=>data_in(65)
   );
   ix25022 : oai21 port map ( Y=>nx25021, A0=>nx36529, A1=>nx42603, B0=>
      nx36531);
   booth_booth_integrtaion_4_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_18, QB=>nx36529, D=>nx25021, CLK=>clk, 
      R=>rst);
   ix36532 : nand03 port map ( Y=>nx36531, A0=>nx42611, A1=>nx9392, A2=>
      nx42607);
   ix9393 : xnor2 port map ( Y=>nx9392, A0=>nx8948, A1=>nx36544);
   ix8949 : oai22 port map ( Y=>nx8948, A0=>nx36514, A1=>nx36535, B0=>
      nx36529, B1=>nx42615);
   ix36538 : aoi32 port map ( Y=>nx36537, A0=>nx8930, A1=>nx41995, A2=>
      nx36540, B0=>data_in(66), B1=>nx41991);
   ix8931 : oai21 port map ( Y=>nx8930, A0=>data_in(64), A1=>data_in(65), B0
      =>data_in(66));
   ix25012 : oai21 port map ( Y=>nx25011, A0=>nx36548, A1=>nx42603, B0=>
      nx36550);
   booth_booth_integrtaion_4_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_19, QB=>nx36548, D=>nx25011, CLK=>clk, 
      R=>rst);
   ix36551 : nand03 port map ( Y=>nx36550, A0=>nx42611, A1=>nx9380, A2=>
      nx42607);
   ix9381 : xnor2 port map ( Y=>nx9380, A0=>nx36553, A1=>nx18382);
   ix36554 : aoi22 port map ( Y=>nx36553, A0=>
      booth_booth_integration_output_4_19, A1=>nx8968, B0=>nx8948, B1=>
      nx18381);
   ix8969 : oai32 port map ( Y=>nx8968, A0=>nx36556, A1=>nx36519, A2=>nx8958, 
      B0=>nx36559, B1=>nx36524);
   ix8935 : nor03_2x port map ( Y=>nx8934, A0=>data_in(66), A1=>data_in(64), 
      A2=>data_in(65));
   ix36560 : inv01 port map ( Y=>nx36559, A=>data_in(67));
   ix8959 : nor04 port map ( Y=>nx8958, A0=>data_in(67), A1=>data_in(66), A2
      =>data_in(64), A3=>data_in(65));
   ix36568 : xnor2 port map ( Y=>nx36567, A0=>nx8996, A1=>nx18383);
   ix8997 : oai22 port map ( Y=>nx8996, A0=>nx36553, A1=>nx36570, B0=>
      nx36581, B1=>nx42617);
   ix36573 : aoi32 port map ( Y=>nx36572, A0=>nx8978, A1=>nx41995, A2=>
      nx36577, B0=>data_in(68), B1=>nx41991);
   ix8979 : nand02 port map ( Y=>nx8978, A0=>nx36575, A1=>data_in(68));
   ix36578 : nand02 port map ( Y=>nx36577, A0=>nx36579, A1=>nx8958);
   ix36580 : inv01 port map ( Y=>nx36579, A=>data_in(68));
   booth_booth_integrtaion_4_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_20, QB=>nx36581, D=>nx25001, CLK=>clk, 
      R=>rst);
   ix24992 : oai21 port map ( Y=>nx24991, A0=>nx36586, A1=>nx42603, B0=>
      nx36588);
   booth_booth_integrtaion_4_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_21, QB=>nx36586, D=>nx24991, CLK=>clk, 
      R=>rst);
   ix36589 : nand03 port map ( Y=>nx36588, A0=>nx42611, A1=>nx9356, A2=>
      nx42607);
   ix9357 : xnor2 port map ( Y=>nx9356, A0=>nx36591, A1=>nx18385);
   ix36592 : aoi22 port map ( Y=>nx36591, A0=>
      booth_booth_integration_output_4_21, A1=>nx9016, B0=>nx8996, B1=>
      nx18383);
   ix9007 : nor02_2x port map ( Y=>nx9006, A0=>data_in(69), A1=>nx36577);
   ix36604 : xnor2 port map ( Y=>nx36603, A0=>nx9044, A1=>nx18386);
   ix9045 : oai22 port map ( Y=>nx9044, A0=>nx36591, A1=>nx36606, B0=>
      nx36617, B1=>nx42619);
   ix36609 : aoi32 port map ( Y=>nx36608, A0=>nx9026, A1=>nx41995, A2=>
      nx36613, B0=>data_in(70), B1=>nx41991);
   ix9027 : nand02 port map ( Y=>nx9026, A0=>nx36611, A1=>data_in(70));
   ix36614 : nand02 port map ( Y=>nx36613, A0=>nx36615, A1=>nx9006);
   ix36616 : inv01 port map ( Y=>nx36615, A=>data_in(70));
   booth_booth_integrtaion_4_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_22, QB=>nx36617, D=>nx24981, CLK=>clk, 
      R=>rst);
   ix24972 : oai21 port map ( Y=>nx24971, A0=>nx36622, A1=>nx42605, B0=>
      nx36624);
   booth_booth_integrtaion_4_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_23, QB=>nx36622, D=>nx24971, CLK=>clk, 
      R=>rst);
   ix36625 : nand03 port map ( Y=>nx36624, A0=>nx42611, A1=>nx9332, A2=>
      nx42607);
   ix9333 : xnor2 port map ( Y=>nx9332, A0=>nx36627, A1=>nx18387);
   ix36628 : aoi22 port map ( Y=>nx36627, A0=>
      booth_booth_integration_output_4_23, A1=>nx9064, B0=>nx9044, B1=>
      nx18386);
   ix9055 : nor02_2x port map ( Y=>nx9054, A0=>data_in(71), A1=>nx36613);
   ix36640 : xnor2 port map ( Y=>nx36639, A0=>nx9092, A1=>nx18388);
   ix9093 : oai22 port map ( Y=>nx9092, A0=>nx36627, A1=>nx36642, B0=>
      nx36653, B1=>nx42621);
   ix36645 : aoi32 port map ( Y=>nx36644, A0=>nx9074, A1=>nx41995, A2=>
      nx36649, B0=>data_in(72), B1=>nx41991);
   ix9075 : nand02 port map ( Y=>nx9074, A0=>nx36647, A1=>data_in(72));
   ix36650 : nand02 port map ( Y=>nx36649, A0=>nx36651, A1=>nx9054);
   ix36652 : inv01 port map ( Y=>nx36651, A=>data_in(72));
   booth_booth_integrtaion_4_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_24, QB=>nx36653, D=>nx24961, CLK=>clk, 
      R=>rst);
   ix24952 : oai21 port map ( Y=>nx24951, A0=>nx36658, A1=>nx42605, B0=>
      nx36660);
   booth_booth_integrtaion_4_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_25, QB=>nx36658, D=>nx24951, CLK=>clk, 
      R=>rst);
   ix36661 : nand03 port map ( Y=>nx36660, A0=>nx42611, A1=>nx9308, A2=>
      nx42607);
   ix9309 : xnor2 port map ( Y=>nx9308, A0=>nx36663, A1=>nx18389);
   ix36664 : aoi22 port map ( Y=>nx36663, A0=>
      booth_booth_integration_output_4_25, A1=>nx9112, B0=>nx9092, B1=>
      nx18388);
   ix9103 : nor02_2x port map ( Y=>nx9102, A0=>data_in(73), A1=>nx36649);
   ix36676 : xnor2 port map ( Y=>nx36675, A0=>nx9140, A1=>nx18390);
   ix9141 : oai22 port map ( Y=>nx9140, A0=>nx36663, A1=>nx36678, B0=>
      nx36689, B1=>nx42623);
   ix36681 : aoi32 port map ( Y=>nx36680, A0=>nx9122, A1=>nx41995, A2=>
      nx36685, B0=>data_in(74), B1=>nx41991);
   ix9123 : nand02 port map ( Y=>nx9122, A0=>nx36683, A1=>data_in(74));
   ix36686 : nand02 port map ( Y=>nx36685, A0=>nx36687, A1=>nx9102);
   ix36688 : inv01 port map ( Y=>nx36687, A=>data_in(74));
   booth_booth_integrtaion_4_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_26, QB=>nx36689, D=>nx24941, CLK=>clk, 
      R=>rst);
   ix24932 : oai21 port map ( Y=>nx24931, A0=>nx36694, A1=>nx42605, B0=>
      nx36696);
   booth_booth_integrtaion_4_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_27, QB=>nx36694, D=>nx24931, CLK=>clk, 
      R=>rst);
   ix36697 : nand03 port map ( Y=>nx36696, A0=>nx43257, A1=>nx9284, A2=>
      nx42607);
   ix9285 : xnor2 port map ( Y=>nx9284, A0=>nx36699, A1=>nx18391);
   ix36700 : aoi22 port map ( Y=>nx36699, A0=>
      booth_booth_integration_output_4_27, A1=>nx9160, B0=>nx9140, B1=>
      nx18390);
   ix9151 : nor02_2x port map ( Y=>nx9150, A0=>data_in(75), A1=>nx36685);
   ix36712 : xnor2 port map ( Y=>nx36711, A0=>nx9188, A1=>nx18393);
   ix9189 : oai22 port map ( Y=>nx9188, A0=>nx36699, A1=>nx36714, B0=>
      nx36725, B1=>nx42625);
   ix36717 : aoi32 port map ( Y=>nx36716, A0=>nx9170, A1=>nx41997, A2=>
      nx36721, B0=>data_in(76), B1=>nx41991);
   ix9171 : nand02 port map ( Y=>nx9170, A0=>nx36719, A1=>data_in(76));
   ix36722 : nand02 port map ( Y=>nx36721, A0=>nx36723, A1=>nx9150);
   ix36724 : inv01 port map ( Y=>nx36723, A=>data_in(76));
   booth_booth_integrtaion_4_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12175, QB=>nx36725, D=>nx24921, CLK=>clk, R=>rst);
   ix24912 : oai21 port map ( Y=>nx24911, A0=>nx36730, A1=>nx42605, B0=>
      nx36732);
   booth_booth_integrtaion_4_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12174, QB=>nx36730, D=>nx24911, CLK=>clk, R=>rst);
   ix36733 : nand03 port map ( Y=>nx36732, A0=>nx43257, A1=>nx9260, A2=>
      nx42605);
   ix9261 : xnor2 port map ( Y=>nx9260, A0=>nx36735, A1=>nx18395);
   ix36736 : aoi22 port map ( Y=>nx36735, A0=>booth_output_29_dup_12174, A1
      =>nx9208, B0=>nx9188, B1=>nx18393);
   ix9199 : nor02_2x port map ( Y=>nx9198, A0=>data_in(77), A1=>nx36721);
   ix24902 : oai21 port map ( Y=>nx24901, A0=>nx36746, A1=>nx42605, B0=>
      nx36748);
   booth_booth_integrtaion_4_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx36746, D=>nx24901, CLK=>clk, R=>rst);
   ix36749 : nand03 port map ( Y=>nx36748, A0=>nx43257, A1=>nx9248, A2=>
      nx42605);
   ix9249 : xnor2 port map ( Y=>nx9248, A0=>nx9236, A1=>nx36763);
   ix9237 : oai22 port map ( Y=>nx9236, A0=>nx36735, A1=>nx36752, B0=>
      nx36746, B1=>nx42627);
   ix36755 : aoi32 port map ( Y=>nx36754, A0=>nx9218, A1=>nx41997, A2=>
      nx36759, B0=>data_in(78), B1=>nx41993);
   ix9219 : nand02 port map ( Y=>nx9218, A0=>nx36757, A1=>data_in(78));
   ix36760 : nand02 port map ( Y=>nx36759, A0=>nx36761, A1=>nx9198);
   ix36762 : inv01 port map ( Y=>nx36761, A=>data_in(78));
   ix9245 : oai22 port map ( Y=>nx9244, A0=>nx36519, A1=>nx36766, B0=>
      nx36768, B1=>nx36524);
   ix36767 : xnor2 port map ( Y=>nx36766, A0=>data_in(79), A1=>nx36759);
   ix36769 : inv01 port map ( Y=>nx36768, A=>data_in(79));
   ix36771 : aoi32 port map ( Y=>nx36770, A0=>nx9194, A1=>nx41997, A2=>
      nx36757, B0=>data_in(77), B1=>nx41993);
   ix9195 : nand02 port map ( Y=>nx9194, A0=>nx36721, A1=>data_in(77));
   ix36774 : aoi32 port map ( Y=>nx36773, A0=>nx9146, A1=>nx41997, A2=>
      nx36719, B0=>data_in(75), B1=>nx41993);
   ix9147 : nand02 port map ( Y=>nx9146, A0=>nx36685, A1=>data_in(75));
   ix36777 : aoi32 port map ( Y=>nx36776, A0=>nx9098, A1=>nx41997, A2=>
      nx36683, B0=>data_in(73), B1=>nx41993);
   ix9099 : nand02 port map ( Y=>nx9098, A0=>nx36649, A1=>data_in(73));
   ix36780 : aoi32 port map ( Y=>nx36779, A0=>nx9050, A1=>nx41997, A2=>
      nx36647, B0=>data_in(71), B1=>nx41993);
   ix9051 : nand02 port map ( Y=>nx9050, A0=>nx36613, A1=>data_in(71));
   ix36783 : aoi32 port map ( Y=>nx36782, A0=>nx9002, A1=>nx41999, A2=>
      nx36611, B0=>data_in(69), B1=>nx41993);
   ix9003 : nand02 port map ( Y=>nx9002, A0=>nx36577, A1=>data_in(69));
   ix36786 : aoi32 port map ( Y=>nx36785, A0=>nx8904, A1=>nx41999, A2=>
      nx36788, B0=>data_in(65), B1=>nx41993);
   ix8905 : nand02 port map ( Y=>nx8904, A0=>data_in(65), A1=>data_in(64));
   booth_booth_integrtaion_4_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_16, QB=>nx36499, D=>nx25041, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_15, QB=>nx36792, D=>nx25051, CLK=>clk, 
      R=>rst);
   ix9485 : aoi21 port map ( Y=>nx9484, A0=>label_5_output_0, A1=>
      booth_booth_integration_output_4_12, B0=>nx43519);
   labelsregfile_label5_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_5_output_1, QB=>nx36809, D=>nx25121, CLK=>clk, R=>rst);
   lat_label_5_input_1 : latch port map ( Q=>label_5_input_1, D=>nx9522, CLK
      =>nx41683);
   reg_label_5_input_state_machine_1 : dffr port map ( Q=>
      label_5_input_state_machine_1, QB=>OPEN, D=>nx25111, CLK=>clk, R=>rst
   );
   ix9519 : xor2 port map ( Y=>nx9518, A0=>nx36350, A1=>nx36799);
   ix36811 : xnor2 port map ( Y=>nx36810, A0=>
      booth_booth_integration_output_4_14, A1=>label_5_output_2);
   labelsregfile_label5_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_5_output_3, QB=>nx36824, D=>nx25161, CLK=>clk, R=>rst);
   lat_label_5_input_3 : latch port map ( Q=>label_5_input_3, D=>nx9586, CLK
      =>nx41683);
   reg_label_5_input_state_machine_3 : dffr port map ( Q=>
      label_5_input_state_machine_3, QB=>OPEN, D=>nx25151, CLK=>clk, R=>rst
   );
   ix9583 : xor2 port map ( Y=>nx9582, A0=>nx36339, A1=>nx36814);
   labelsregfile_label5_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_5_output_5, QB=>nx36839, D=>nx25201, CLK=>clk, R=>rst);
   lat_label_5_input_5 : latch port map ( Q=>label_5_input_5, D=>nx9650, CLK
      =>nx41683);
   reg_label_5_input_state_machine_5 : dffr port map ( Q=>
      label_5_input_state_machine_5, QB=>OPEN, D=>nx25191, CLK=>clk, R=>rst
   );
   ix9647 : xor2 port map ( Y=>nx9646, A0=>nx36328, A1=>nx36829);
   labelsregfile_label5_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_5_output_7, QB=>nx36854, D=>nx25241, CLK=>clk, R=>rst);
   lat_label_5_input_7 : latch port map ( Q=>label_5_input_7, D=>nx9714, CLK
      =>nx41685);
   reg_label_5_input_state_machine_7 : dffr port map ( Q=>
      label_5_input_state_machine_7, QB=>OPEN, D=>nx25231, CLK=>clk, R=>rst
   );
   ix9711 : xor2 port map ( Y=>nx9710, A0=>nx36317, A1=>nx36844);
   labelsregfile_label5_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_5_output_9, QB=>nx36869, D=>nx25281, CLK=>clk, R=>rst);
   lat_label_5_input_9 : latch port map ( Q=>label_5_input_9, D=>nx9778, CLK
      =>nx41685);
   reg_label_5_input_state_machine_9 : dffr port map ( Q=>
      label_5_input_state_machine_9, QB=>OPEN, D=>nx25271, CLK=>clk, R=>rst
   );
   ix9775 : xor2 port map ( Y=>nx9774, A0=>nx36306, A1=>nx36859);
   labelsregfile_label5_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_5_output_11, QB=>nx36884, D=>nx25321, CLK=>clk, R=>rst);
   lat_label_5_input_11 : latch port map ( Q=>label_5_input_11, D=>nx9842, 
      CLK=>nx41685);
   reg_label_5_input_state_machine_11 : dffr port map ( Q=>
      label_5_input_state_machine_11, QB=>OPEN, D=>nx25311, CLK=>clk, R=>rst
   );
   ix9839 : xor2 port map ( Y=>nx9838, A0=>nx36295, A1=>nx36874);
   labelsregfile_label5_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_5_output_13, QB=>nx36899, D=>nx25361, CLK=>clk, R=>rst);
   lat_label_5_input_13 : latch port map ( Q=>label_5_input_13, D=>nx9906, 
      CLK=>nx41687);
   reg_label_5_input_state_machine_13 : dffr port map ( Q=>
      label_5_input_state_machine_13, QB=>OPEN, D=>nx25351, CLK=>clk, R=>rst
   );
   ix9903 : xor2 port map ( Y=>nx9902, A0=>nx36284, A1=>nx36889);
   ix36904 : nor03_2x port map ( Y=>nx36903, A0=>nx41565, A1=>nx41371, A2=>
      nx1782);
   ix26222 : oai21 port map ( Y=>nx26221, A0=>nx36907, A1=>nx41605, B0=>
      nx36909);
   max_calc_reg_comparator_third_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx36907, D=>nx26221, CLK=>clk);
   ix36910 : nand03 port map ( Y=>nx36909, A0=>label_6_output_14, A1=>
      nx42631, A2=>nx41605);
   labelsregfile_label6_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_6_output_14, QB=>OPEN, D=>nx26211, CLK=>clk, R=>rst);
   lat_label_6_input_14 : latch port map ( Q=>label_6_input_14, D=>nx11250, 
      CLK=>nx41691);
   reg_label_6_input_state_machine_14 : dffr port map ( Q=>
      label_6_input_state_machine_14, QB=>OPEN, D=>nx25391, CLK=>clk, R=>rst
   );
   ix11247 : xnor2 port map ( Y=>nx11246, A0=>nx11242, A1=>nx37536);
   ix11243 : oai22 port map ( Y=>nx11242, A0=>nx36920, A1=>nx37525, B0=>
      nx37535, B1=>nx37294);
   ix36921 : aoi22 port map ( Y=>nx36920, A0=>label_6_output_12, A1=>
      booth_booth_integration_output_5_24, B0=>nx11178, B1=>nx18457);
   labelsregfile_label6_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_6_output_12, QB=>OPEN, D=>nx26181, CLK=>clk, R=>rst);
   lat_label_6_input_12 : latch port map ( Q=>label_6_input_12, D=>nx11192, 
      CLK=>nx41691);
   reg_label_6_input_state_machine_12 : dffr port map ( Q=>
      label_6_input_state_machine_12, QB=>OPEN, D=>nx26171, CLK=>clk, R=>rst
   );
   ix11189 : xnor2 port map ( Y=>nx11188, A0=>nx11178, A1=>nx37521);
   ix11179 : oai22 port map ( Y=>nx11178, A0=>nx36931, A1=>nx37510, B0=>
      nx37520, B1=>nx37258);
   ix36932 : aoi22 port map ( Y=>nx36931, A0=>label_6_output_10, A1=>
      booth_booth_integration_output_5_22, B0=>nx11114, B1=>nx18455);
   labelsregfile_label6_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_6_output_10, QB=>OPEN, D=>nx26141, CLK=>clk, R=>rst);
   lat_label_6_input_10 : latch port map ( Q=>label_6_input_10, D=>nx11128, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_10 : dffr port map ( Q=>
      label_6_input_state_machine_10, QB=>OPEN, D=>nx26131, CLK=>clk, R=>rst
   );
   ix11125 : xnor2 port map ( Y=>nx11124, A0=>nx11114, A1=>nx37506);
   ix11115 : oai22 port map ( Y=>nx11114, A0=>nx36942, A1=>nx37495, B0=>
      nx37505, B1=>nx37222);
   ix36943 : aoi22 port map ( Y=>nx36942, A0=>label_6_output_8, A1=>
      booth_booth_integration_output_5_20, B0=>nx11050, B1=>nx18453);
   labelsregfile_label6_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_6_output_8, QB=>OPEN, D=>nx26101, CLK=>clk, R=>rst);
   lat_label_6_input_8 : latch port map ( Q=>label_6_input_8, D=>nx11064, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_8 : dffr port map ( Q=>
      label_6_input_state_machine_8, QB=>OPEN, D=>nx26091, CLK=>clk, R=>rst
   );
   ix11061 : xnor2 port map ( Y=>nx11060, A0=>nx11050, A1=>nx37491);
   ix11051 : oai22 port map ( Y=>nx11050, A0=>nx36953, A1=>nx37480, B0=>
      nx37490, B1=>nx37184);
   ix36954 : aoi22 port map ( Y=>nx36953, A0=>label_6_output_6, A1=>
      booth_booth_integration_output_5_18, B0=>nx10986, B1=>nx18449);
   labelsregfile_label6_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_6_output_6, QB=>OPEN, D=>nx26061, CLK=>clk, R=>rst);
   lat_label_6_input_6 : latch port map ( Q=>label_6_input_6, D=>nx11000, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_6 : dffr port map ( Q=>
      label_6_input_state_machine_6, QB=>OPEN, D=>nx26051, CLK=>clk, R=>rst
   );
   ix10997 : xnor2 port map ( Y=>nx10996, A0=>nx10986, A1=>nx37476);
   ix10987 : oai22 port map ( Y=>nx10986, A0=>nx36964, A1=>nx37465, B0=>
      nx37475, B1=>nx37145);
   ix36965 : aoi22 port map ( Y=>nx36964, A0=>label_6_output_4, A1=>
      booth_booth_integration_output_5_16, B0=>nx10922, B1=>nx18445);
   labelsregfile_label6_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_6_output_4, QB=>OPEN, D=>nx26021, CLK=>clk, R=>rst);
   lat_label_6_input_4 : latch port map ( Q=>label_6_input_4, D=>nx10936, 
      CLK=>nx41687);
   reg_label_6_input_state_machine_4 : dffr port map ( Q=>
      label_6_input_state_machine_4, QB=>OPEN, D=>nx26011, CLK=>clk, R=>rst
   );
   ix10933 : xnor2 port map ( Y=>nx10932, A0=>nx10922, A1=>nx37461);
   ix10923 : oai22 port map ( Y=>nx10922, A0=>nx36975, A1=>nx37450, B0=>
      nx37460, B1=>nx37428);
   ix36976 : aoi22 port map ( Y=>nx36975, A0=>label_6_output_2, A1=>
      booth_booth_integration_output_5_14, B0=>nx10858, B1=>nx18443);
   labelsregfile_label6_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_6_output_2, QB=>OPEN, D=>nx25981, CLK=>clk, R=>rst);
   lat_label_6_input_2 : latch port map ( Q=>label_6_input_2, D=>nx10872, 
      CLK=>nx41687);
   reg_label_6_input_state_machine_2 : dffr port map ( Q=>
      label_6_input_state_machine_2, QB=>OPEN, D=>nx25971, CLK=>clk, R=>rst
   );
   ix10869 : xnor2 port map ( Y=>nx10868, A0=>nx10858, A1=>nx37446);
   ix10859 : oai22 port map ( Y=>nx10858, A0=>nx36986, A1=>nx37435, B0=>
      nx37445, B1=>nx37431);
   ix36987 : nand02 port map ( Y=>nx36986, A0=>label_6_output_0, A1=>
      booth_booth_integration_output_5_12);
   labelsregfile_label6_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_6_output_0, QB=>OPEN, D=>nx25941, CLK=>clk, R=>rst);
   lat_label_6_input_0 : latch port map ( Q=>label_6_input_0, D=>nx10814, 
      CLK=>nx41687);
   ix10815 : oai21 port map ( Y=>nx10814, A0=>nx36992, A1=>nx41447, B0=>
      nx36996);
   reg_label_6_input_state_machine_0 : dffr port map ( Q=>
      label_6_input_state_machine_0, QB=>nx36992, D=>nx25931, CLK=>clk, R=>
      rst);
   ix36997 : oai21 port map ( Y=>nx36996, A0=>
      booth_booth_integration_output_5_12, A1=>label_6_output_0, B0=>nx10802
   );
   booth_booth_integrtaion_5_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_12, QB=>OPEN, D=>nx25921, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_13, QB=>nx37431, D=>nx25911, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_14, QB=>OPEN, D=>nx25901, CLK=>clk, R
      =>rst);
   ix37010 : aoi22 port map ( Y=>nx37009, A0=>nx41797, A1=>nx42015, B0=>
      nx10744, B1=>nx10750);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_reg_output_0, QB=>OPEN, 
      D=>nx25421, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_0, QB=>OPEN, D=>nx25407, CLK
      =>clk, S=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_reg_output_9, QB=>OPEN, 
      D=>nx25601, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_9, QB=>OPEN, D=>nx25591, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12828, QB=>OPEN, D=>nx25581, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_8, QB=>OPEN, D=>nx25571, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12829, QB=>OPEN, D=>nx25561, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_7, QB=>OPEN, D=>nx25551, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12830, QB=>OPEN, D=>nx25541, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_6, QB=>OPEN, D=>nx25531, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12831, QB=>OPEN, D=>nx25521, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_5, QB=>OPEN, D=>nx25511, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12832, QB=>OPEN, D=>nx25501, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_4, QB=>OPEN, D=>nx25491, CLK
      =>clk, R=>nx41495);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12833, QB=>OPEN, D=>nx25481, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_3, QB=>OPEN, D=>nx25471, CLK
      =>clk, R=>nx41493);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12834, QB=>OPEN, D=>nx25461, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_2, QB=>OPEN, D=>nx25451, CLK
      =>clk, R=>nx41493);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12835, QB=>OPEN, D=>nx25441, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_1, QB=>OPEN, D=>nx25431, CLK
      =>clk, R=>nx41493);
   ix25402 : nand02 port map ( Y=>nx25401, A0=>nx42949, A1=>nx42001);
   booth_booth_integrtaion_5_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx37056, D=>nx25401, CLK=>clk, S=>nx41493);
   ix10745 : nand02 port map ( Y=>nx10744, A0=>nx37077, A1=>nx37135);
   ix37078 : oai21 port map ( Y=>nx37077, A0=>nx42027, A1=>nx42023, B0=>
      data_in(80));
   ix25732 : oai21 port map ( Y=>nx25731, A0=>nx37082, A1=>nx42651, B0=>
      nx37084);
   booth_booth_integrtaion_5_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx37082, D=>nx25731, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12206, QB=>nx37133, D=>nx25721, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12205, QB=>OPEN, D=>nx25711, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12204, QB=>OPEN, D=>nx25701, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12203, QB=>OPEN, D=>nx25691, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12202, QB=>OPEN, D=>nx25681, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12201, QB=>OPEN, D=>nx25671, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12200, QB=>OPEN, D=>nx25661, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12199, QB=>OPEN, D=>nx25651, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12198, QB=>OPEN, D=>nx25641, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12197, QB=>OPEN, D=>nx25631, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12196, QB=>OPEN, D=>nx25621, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12195, QB=>OPEN, D=>nx25611, CLK=>clk, R=>rst);
   ix37140 : xnor2 port map ( Y=>nx37139, A0=>nx10214, A1=>nx18421);
   ix25872 : oai21 port map ( Y=>nx25871, A0=>nx37145, A1=>nx42651, B0=>
      nx37147);
   booth_booth_integrtaion_5_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_17, QB=>nx37145, D=>nx25871, CLK=>clk, 
      R=>rst);
   ix37148 : nand03 port map ( Y=>nx37147, A0=>nx42659, A1=>nx10722, A2=>
      nx42655);
   ix10723 : xnor2 port map ( Y=>nx10722, A0=>nx37150, A1=>nx18422);
   ix37151 : aoi22 port map ( Y=>nx37150, A0=>
      booth_booth_integration_output_5_17, A1=>nx10238, B0=>nx10214, B1=>
      nx18421);
   ix10229 : nor02_2x port map ( Y=>nx10228, A0=>data_in(80), A1=>
      data_in(81));
   ix25862 : oai21 port map ( Y=>nx25861, A0=>nx37165, A1=>nx42651, B0=>
      nx37167);
   booth_booth_integrtaion_5_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_18, QB=>nx37165, D=>nx25861, CLK=>clk, 
      R=>rst);
   ix37168 : nand03 port map ( Y=>nx37167, A0=>nx42659, A1=>nx10710, A2=>
      nx42655);
   ix10711 : xnor2 port map ( Y=>nx10710, A0=>nx10266, A1=>nx37180);
   ix10267 : oai22 port map ( Y=>nx10266, A0=>nx37150, A1=>nx37171, B0=>
      nx37165, B1=>nx42663);
   ix37174 : aoi32 port map ( Y=>nx37173, A0=>nx10248, A1=>nx42027, A2=>
      nx37176, B0=>data_in(82), B1=>nx42023);
   ix10249 : oai21 port map ( Y=>nx10248, A0=>data_in(80), A1=>data_in(81), 
      B0=>data_in(82));
   ix25852 : oai21 port map ( Y=>nx25851, A0=>nx37184, A1=>nx42651, B0=>
      nx37186);
   booth_booth_integrtaion_5_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_19, QB=>nx37184, D=>nx25851, CLK=>clk, 
      R=>rst);
   ix37187 : nand03 port map ( Y=>nx37186, A0=>nx42659, A1=>nx10698, A2=>
      nx42655);
   ix10699 : xnor2 port map ( Y=>nx10698, A0=>nx37189, A1=>nx18424);
   ix37190 : aoi22 port map ( Y=>nx37189, A0=>
      booth_booth_integration_output_5_19, A1=>nx10286, B0=>nx10266, B1=>
      nx18423);
   ix10287 : oai32 port map ( Y=>nx10286, A0=>nx37192, A1=>nx37155, A2=>
      nx10276, B0=>nx37195, B1=>nx37160);
   ix10253 : nor03_2x port map ( Y=>nx10252, A0=>data_in(82), A1=>
      data_in(80), A2=>data_in(81));
   ix37196 : inv01 port map ( Y=>nx37195, A=>data_in(83));
   ix10277 : nor04 port map ( Y=>nx10276, A0=>data_in(83), A1=>data_in(82), 
      A2=>data_in(80), A3=>data_in(81));
   ix37204 : xnor2 port map ( Y=>nx37203, A0=>nx10314, A1=>nx18425);
   ix10315 : oai22 port map ( Y=>nx10314, A0=>nx37189, A1=>nx37206, B0=>
      nx37217, B1=>nx42665);
   ix37209 : aoi32 port map ( Y=>nx37208, A0=>nx10296, A1=>nx42027, A2=>
      nx37213, B0=>data_in(84), B1=>nx42023);
   ix10297 : nand02 port map ( Y=>nx10296, A0=>nx37211, A1=>data_in(84));
   ix37214 : nand02 port map ( Y=>nx37213, A0=>nx37215, A1=>nx10276);
   ix37216 : inv01 port map ( Y=>nx37215, A=>data_in(84));
   booth_booth_integrtaion_5_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_20, QB=>nx37217, D=>nx25841, CLK=>clk, 
      R=>rst);
   ix25832 : oai21 port map ( Y=>nx25831, A0=>nx37222, A1=>nx42651, B0=>
      nx37224);
   booth_booth_integrtaion_5_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_21, QB=>nx37222, D=>nx25831, CLK=>clk, 
      R=>rst);
   ix37225 : nand03 port map ( Y=>nx37224, A0=>nx42659, A1=>nx10674, A2=>
      nx42655);
   ix10675 : xnor2 port map ( Y=>nx10674, A0=>nx37227, A1=>nx18426);
   ix37228 : aoi22 port map ( Y=>nx37227, A0=>
      booth_booth_integration_output_5_21, A1=>nx10334, B0=>nx10314, B1=>
      nx18425);
   ix10325 : nor02_2x port map ( Y=>nx10324, A0=>data_in(85), A1=>nx37213);
   ix37240 : xnor2 port map ( Y=>nx37239, A0=>nx10362, A1=>nx18427);
   ix10363 : oai22 port map ( Y=>nx10362, A0=>nx37227, A1=>nx37242, B0=>
      nx37253, B1=>nx42667);
   ix37245 : aoi32 port map ( Y=>nx37244, A0=>nx10344, A1=>nx42027, A2=>
      nx37249, B0=>data_in(86), B1=>nx42023);
   ix10345 : nand02 port map ( Y=>nx10344, A0=>nx37247, A1=>data_in(86));
   ix37250 : nand02 port map ( Y=>nx37249, A0=>nx37251, A1=>nx10324);
   ix37252 : inv01 port map ( Y=>nx37251, A=>data_in(86));
   booth_booth_integrtaion_5_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_22, QB=>nx37253, D=>nx25821, CLK=>clk, 
      R=>rst);
   ix25812 : oai21 port map ( Y=>nx25811, A0=>nx37258, A1=>nx42653, B0=>
      nx37260);
   booth_booth_integrtaion_5_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_23, QB=>nx37258, D=>nx25811, CLK=>clk, 
      R=>rst);
   ix37261 : nand03 port map ( Y=>nx37260, A0=>nx42659, A1=>nx10650, A2=>
      nx42655);
   ix10651 : xnor2 port map ( Y=>nx10650, A0=>nx37263, A1=>nx18429);
   ix37264 : aoi22 port map ( Y=>nx37263, A0=>
      booth_booth_integration_output_5_23, A1=>nx10382, B0=>nx10362, B1=>
      nx18427);
   ix10373 : nor02_2x port map ( Y=>nx10372, A0=>data_in(87), A1=>nx37249);
   ix37276 : xnor2 port map ( Y=>nx37275, A0=>nx10410, A1=>nx18431);
   ix10411 : oai22 port map ( Y=>nx10410, A0=>nx37263, A1=>nx37278, B0=>
      nx37289, B1=>nx42669);
   ix37281 : aoi32 port map ( Y=>nx37280, A0=>nx10392, A1=>nx42027, A2=>
      nx37285, B0=>data_in(88), B1=>nx42023);
   ix10393 : nand02 port map ( Y=>nx10392, A0=>nx37283, A1=>data_in(88));
   ix37286 : nand02 port map ( Y=>nx37285, A0=>nx37287, A1=>nx10372);
   ix37288 : inv01 port map ( Y=>nx37287, A=>data_in(88));
   booth_booth_integrtaion_5_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_24, QB=>nx37289, D=>nx25801, CLK=>clk, 
      R=>rst);
   ix25792 : oai21 port map ( Y=>nx25791, A0=>nx37294, A1=>nx42653, B0=>
      nx37296);
   booth_booth_integrtaion_5_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_25, QB=>nx37294, D=>nx25791, CLK=>clk, 
      R=>rst);
   ix37297 : nand03 port map ( Y=>nx37296, A0=>nx42659, A1=>nx10626, A2=>
      nx42655);
   ix10627 : xnor2 port map ( Y=>nx10626, A0=>nx37299, A1=>nx18433);
   ix37300 : aoi22 port map ( Y=>nx37299, A0=>
      booth_booth_integration_output_5_25, A1=>nx10430, B0=>nx10410, B1=>
      nx18431);
   ix10421 : nor02_2x port map ( Y=>nx10420, A0=>data_in(89), A1=>nx37285);
   ix37312 : xnor2 port map ( Y=>nx37311, A0=>nx10458, A1=>nx18435);
   ix10459 : oai22 port map ( Y=>nx10458, A0=>nx37299, A1=>nx37314, B0=>
      nx37325, B1=>nx42671);
   ix37317 : aoi32 port map ( Y=>nx37316, A0=>nx10440, A1=>nx42027, A2=>
      nx37321, B0=>data_in(90), B1=>nx42023);
   ix10441 : nand02 port map ( Y=>nx10440, A0=>nx37319, A1=>data_in(90));
   ix37322 : nand02 port map ( Y=>nx37321, A0=>nx37323, A1=>nx10420);
   ix37324 : inv01 port map ( Y=>nx37323, A=>data_in(90));
   booth_booth_integrtaion_5_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_26, QB=>nx37325, D=>nx25781, CLK=>clk, 
      R=>rst);
   ix25772 : oai21 port map ( Y=>nx25771, A0=>nx37330, A1=>nx42653, B0=>
      nx37332);
   booth_booth_integrtaion_5_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_27, QB=>nx37330, D=>nx25771, CLK=>clk, 
      R=>rst);
   ix37333 : nand03 port map ( Y=>nx37332, A0=>nx43277, A1=>nx10602, A2=>
      nx42655);
   ix10603 : xnor2 port map ( Y=>nx10602, A0=>nx37335, A1=>nx18437);
   ix37336 : aoi22 port map ( Y=>nx37335, A0=>
      booth_booth_integration_output_5_27, A1=>nx10478, B0=>nx10458, B1=>
      nx18435);
   ix10469 : nor02_2x port map ( Y=>nx10468, A0=>data_in(91), A1=>nx37321);
   ix37348 : xnor2 port map ( Y=>nx37347, A0=>nx10506, A1=>nx18439);
   ix10507 : oai22 port map ( Y=>nx10506, A0=>nx37335, A1=>nx37350, B0=>
      nx37361, B1=>nx42673);
   ix37353 : aoi32 port map ( Y=>nx37352, A0=>nx10488, A1=>nx42029, A2=>
      nx37357, B0=>data_in(92), B1=>nx42023);
   ix10489 : nand02 port map ( Y=>nx10488, A0=>nx37355, A1=>data_in(92));
   ix37358 : nand02 port map ( Y=>nx37357, A0=>nx37359, A1=>nx10468);
   ix37360 : inv01 port map ( Y=>nx37359, A=>data_in(92));
   booth_booth_integrtaion_5_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12194, QB=>nx37361, D=>nx25761, CLK=>clk, R=>rst);
   ix25752 : oai21 port map ( Y=>nx25751, A0=>nx37366, A1=>nx42653, B0=>
      nx37368);
   booth_booth_integrtaion_5_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12193, QB=>nx37366, D=>nx25751, CLK=>clk, R=>rst);
   ix37369 : nand03 port map ( Y=>nx37368, A0=>nx43277, A1=>nx10578, A2=>
      nx42653);
   ix10579 : xnor2 port map ( Y=>nx10578, A0=>nx37371, A1=>nx18440);
   ix37372 : aoi22 port map ( Y=>nx37371, A0=>booth_output_29_dup_12193, A1
      =>nx10526, B0=>nx10506, B1=>nx18439);
   ix10517 : nor02_2x port map ( Y=>nx10516, A0=>data_in(93), A1=>nx37357);
   ix25742 : oai21 port map ( Y=>nx25741, A0=>nx37382, A1=>nx42653, B0=>
      nx37384);
   booth_booth_integrtaion_5_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx37382, D=>nx25741, CLK=>clk, R=>rst);
   ix37385 : nand03 port map ( Y=>nx37384, A0=>nx43277, A1=>nx10566, A2=>
      nx42653);
   ix10567 : xnor2 port map ( Y=>nx10566, A0=>nx10554, A1=>nx37399);
   ix10555 : oai22 port map ( Y=>nx10554, A0=>nx37371, A1=>nx37388, B0=>
      nx37382, B1=>nx42675);
   ix37391 : aoi32 port map ( Y=>nx37390, A0=>nx10536, A1=>nx42029, A2=>
      nx37395, B0=>data_in(94), B1=>nx42025);
   ix10537 : nand02 port map ( Y=>nx10536, A0=>nx37393, A1=>data_in(94));
   ix37396 : nand02 port map ( Y=>nx37395, A0=>nx37397, A1=>nx10516);
   ix37398 : inv01 port map ( Y=>nx37397, A=>data_in(94));
   ix10563 : oai22 port map ( Y=>nx10562, A0=>nx37155, A1=>nx37402, B0=>
      nx37404, B1=>nx37160);
   ix37403 : xnor2 port map ( Y=>nx37402, A0=>data_in(95), A1=>nx37395);
   ix37405 : inv01 port map ( Y=>nx37404, A=>data_in(95));
   ix37407 : aoi32 port map ( Y=>nx37406, A0=>nx10512, A1=>nx42029, A2=>
      nx37393, B0=>data_in(93), B1=>nx42025);
   ix10513 : nand02 port map ( Y=>nx10512, A0=>nx37357, A1=>data_in(93));
   ix37410 : aoi32 port map ( Y=>nx37409, A0=>nx10464, A1=>nx42029, A2=>
      nx37355, B0=>data_in(91), B1=>nx42025);
   ix10465 : nand02 port map ( Y=>nx10464, A0=>nx37321, A1=>data_in(91));
   ix37413 : aoi32 port map ( Y=>nx37412, A0=>nx10416, A1=>nx42029, A2=>
      nx37319, B0=>data_in(89), B1=>nx42025);
   ix10417 : nand02 port map ( Y=>nx10416, A0=>nx37285, A1=>data_in(89));
   ix37416 : aoi32 port map ( Y=>nx37415, A0=>nx10368, A1=>nx42029, A2=>
      nx37283, B0=>data_in(87), B1=>nx42025);
   ix10369 : nand02 port map ( Y=>nx10368, A0=>nx37249, A1=>data_in(87));
   ix37419 : aoi32 port map ( Y=>nx37418, A0=>nx10320, A1=>nx42031, A2=>
      nx37247, B0=>data_in(85), B1=>nx42025);
   ix10321 : nand02 port map ( Y=>nx10320, A0=>nx37213, A1=>data_in(85));
   ix37422 : aoi32 port map ( Y=>nx37421, A0=>nx10222, A1=>nx42031, A2=>
      nx37424, B0=>data_in(81), B1=>nx42025);
   ix10223 : nand02 port map ( Y=>nx10222, A0=>data_in(81), A1=>data_in(80)
   );
   booth_booth_integrtaion_5_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_16, QB=>nx37135, D=>nx25881, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_15, QB=>nx37428, D=>nx25891, CLK=>clk, 
      R=>rst);
   ix10803 : aoi21 port map ( Y=>nx10802, A0=>label_6_output_0, A1=>
      booth_booth_integration_output_5_12, B0=>nx43055);
   labelsregfile_label6_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_6_output_1, QB=>nx37445, D=>nx25961, CLK=>clk, R=>rst);
   lat_label_6_input_1 : latch port map ( Q=>label_6_input_1, D=>nx10840, 
      CLK=>nx41687);
   reg_label_6_input_state_machine_1 : dffr port map ( Q=>
      label_6_input_state_machine_1, QB=>OPEN, D=>nx25951, CLK=>clk, R=>rst
   );
   ix10837 : xor2 port map ( Y=>nx10836, A0=>nx36986, A1=>nx37435);
   ix37447 : xnor2 port map ( Y=>nx37446, A0=>
      booth_booth_integration_output_5_14, A1=>label_6_output_2);
   labelsregfile_label6_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_6_output_3, QB=>nx37460, D=>nx26001, CLK=>clk, R=>rst);
   lat_label_6_input_3 : latch port map ( Q=>label_6_input_3, D=>nx10904, 
      CLK=>nx41687);
   reg_label_6_input_state_machine_3 : dffr port map ( Q=>
      label_6_input_state_machine_3, QB=>OPEN, D=>nx25991, CLK=>clk, R=>rst
   );
   ix10901 : xor2 port map ( Y=>nx10900, A0=>nx36975, A1=>nx37450);
   labelsregfile_label6_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_6_output_5, QB=>nx37475, D=>nx26041, CLK=>clk, R=>rst);
   lat_label_6_input_5 : latch port map ( Q=>label_6_input_5, D=>nx10968, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_5 : dffr port map ( Q=>
      label_6_input_state_machine_5, QB=>OPEN, D=>nx26031, CLK=>clk, R=>rst
   );
   ix10965 : xor2 port map ( Y=>nx10964, A0=>nx36964, A1=>nx37465);
   labelsregfile_label6_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_6_output_7, QB=>nx37490, D=>nx26081, CLK=>clk, R=>rst);
   lat_label_6_input_7 : latch port map ( Q=>label_6_input_7, D=>nx11032, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_7 : dffr port map ( Q=>
      label_6_input_state_machine_7, QB=>OPEN, D=>nx26071, CLK=>clk, R=>rst
   );
   ix11029 : xor2 port map ( Y=>nx11028, A0=>nx36953, A1=>nx37480);
   labelsregfile_label6_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_6_output_9, QB=>nx37505, D=>nx26121, CLK=>clk, R=>rst);
   lat_label_6_input_9 : latch port map ( Q=>label_6_input_9, D=>nx11096, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_9 : dffr port map ( Q=>
      label_6_input_state_machine_9, QB=>OPEN, D=>nx26111, CLK=>clk, R=>rst
   );
   ix11093 : xor2 port map ( Y=>nx11092, A0=>nx36942, A1=>nx37495);
   labelsregfile_label6_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_6_output_11, QB=>nx37520, D=>nx26161, CLK=>clk, R=>rst);
   lat_label_6_input_11 : latch port map ( Q=>label_6_input_11, D=>nx11160, 
      CLK=>nx41689);
   reg_label_6_input_state_machine_11 : dffr port map ( Q=>
      label_6_input_state_machine_11, QB=>OPEN, D=>nx26151, CLK=>clk, R=>rst
   );
   ix11157 : xor2 port map ( Y=>nx11156, A0=>nx36931, A1=>nx37510);
   labelsregfile_label6_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_6_output_13, QB=>nx37535, D=>nx26201, CLK=>clk, R=>rst);
   lat_label_6_input_13 : latch port map ( Q=>label_6_input_13, D=>nx11224, 
      CLK=>nx41691);
   reg_label_6_input_state_machine_13 : dffr port map ( Q=>
      label_6_input_state_machine_13, QB=>OPEN, D=>nx26191, CLK=>clk, R=>rst
   );
   ix11221 : xor2 port map ( Y=>nx11220, A0=>nx36920, A1=>nx37525);
   ix11787 : xnor2 port map ( Y=>nx11786, A0=>nx37540, A1=>nx11784);
   ix37541 : aoi22 port map ( Y=>nx37540, A0=>nx36907, A1=>
      max_calc_comparator_third_inp1_14, B0=>nx11272, B1=>nx11690);
   ix11691 : oai22 port map ( Y=>nx11690, A0=>nx37544, A1=>nx37557, B0=>
      max_calc_comparator_third_inp2_13, B1=>nx37552);
   ix26232 : oai21 port map ( Y=>nx26231, A0=>nx37548, A1=>nx41605, B0=>
      nx37550);
   max_calc_reg_comparator_third_inp2_13 : dff port map ( Q=>
      max_calc_comparator_third_inp2_13, QB=>nx37548, D=>nx26231, CLK=>clk);
   max_calc_reg_comparator_third_inp1_13 : dff port map ( Q=>
      max_calc_comparator_third_inp1_13, QB=>nx37552, D=>nx26241, CLK=>clk);
   ix26242 : oai21 port map ( Y=>nx26241, A0=>nx37552, A1=>nx41607, B0=>
      nx37555);
   ix37558 : aoi22 port map ( Y=>nx37557, A0=>nx37559, A1=>
      max_calc_comparator_third_inp1_12, B0=>nx11316, B1=>nx11674);
   max_calc_reg_comparator_third_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx37559, D=>nx26251, CLK=>clk);
   ix26252 : oai21 port map ( Y=>nx26251, A0=>nx37559, A1=>nx41607, B0=>
      nx37562);
   ix37563 : nand03 port map ( Y=>nx37562, A0=>label_6_output_12, A1=>
      nx42631, A2=>nx41607);
   ix26262 : oai21 port map ( Y=>nx26261, A0=>nx37566, A1=>nx41607, B0=>
      nx37568);
   max_calc_reg_comparator_third_inp1_12 : dff port map ( Q=>
      max_calc_comparator_third_inp1_12, QB=>nx37566, D=>nx26261, CLK=>clk);
   ix37569 : nand03 port map ( Y=>nx37568, A0=>label_5_output_12, A1=>
      nx42631, A2=>nx41607);
   ix11675 : oai22 port map ( Y=>nx11674, A0=>nx37572, A1=>nx37585, B0=>
      max_calc_comparator_third_inp2_11, B1=>nx37580);
   ix26272 : oai21 port map ( Y=>nx26271, A0=>nx37576, A1=>nx41609, B0=>
      nx37578);
   max_calc_reg_comparator_third_inp2_11 : dff port map ( Q=>
      max_calc_comparator_third_inp2_11, QB=>nx37576, D=>nx26271, CLK=>clk);
   max_calc_reg_comparator_third_inp1_11 : dff port map ( Q=>
      max_calc_comparator_third_inp1_11, QB=>nx37580, D=>nx26281, CLK=>clk);
   ix26282 : oai21 port map ( Y=>nx26281, A0=>nx37580, A1=>nx41609, B0=>
      nx37583);
   ix37586 : aoi22 port map ( Y=>nx37585, A0=>nx37587, A1=>
      max_calc_comparator_third_inp1_10, B0=>nx11360, B1=>nx11658);
   max_calc_reg_comparator_third_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx37587, D=>nx26291, CLK=>clk);
   ix26292 : oai21 port map ( Y=>nx26291, A0=>nx37587, A1=>nx41609, B0=>
      nx37590);
   ix37591 : nand03 port map ( Y=>nx37590, A0=>label_6_output_10, A1=>
      nx42633, A2=>nx41609);
   ix26302 : oai21 port map ( Y=>nx26301, A0=>nx37594, A1=>nx41609, B0=>
      nx37596);
   max_calc_reg_comparator_third_inp1_10 : dff port map ( Q=>
      max_calc_comparator_third_inp1_10, QB=>nx37594, D=>nx26301, CLK=>clk);
   ix37597 : nand03 port map ( Y=>nx37596, A0=>label_5_output_10, A1=>
      nx42633, A2=>nx41611);
   ix11659 : oai22 port map ( Y=>nx11658, A0=>nx37600, A1=>nx37613, B0=>
      max_calc_comparator_third_inp2_9, B1=>nx37608);
   ix26312 : oai21 port map ( Y=>nx26311, A0=>nx37604, A1=>nx41611, B0=>
      nx37606);
   max_calc_reg_comparator_third_inp2_9 : dff port map ( Q=>
      max_calc_comparator_third_inp2_9, QB=>nx37604, D=>nx26311, CLK=>clk);
   max_calc_reg_comparator_third_inp1_9 : dff port map ( Q=>
      max_calc_comparator_third_inp1_9, QB=>nx37608, D=>nx26321, CLK=>clk);
   ix26322 : oai21 port map ( Y=>nx26321, A0=>nx37608, A1=>nx41611, B0=>
      nx37611);
   ix37614 : aoi22 port map ( Y=>nx37613, A0=>nx37615, A1=>
      max_calc_comparator_third_inp1_8, B0=>nx11404, B1=>nx11642);
   max_calc_reg_comparator_third_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx37615, D=>nx26331, CLK=>clk);
   ix26332 : oai21 port map ( Y=>nx26331, A0=>nx37615, A1=>nx41611, B0=>
      nx37618);
   ix37619 : nand03 port map ( Y=>nx37618, A0=>label_6_output_8, A1=>nx42633, 
      A2=>nx41611);
   ix26342 : oai21 port map ( Y=>nx26341, A0=>nx37622, A1=>nx41613, B0=>
      nx37624);
   max_calc_reg_comparator_third_inp1_8 : dff port map ( Q=>
      max_calc_comparator_third_inp1_8, QB=>nx37622, D=>nx26341, CLK=>clk);
   ix37625 : nand03 port map ( Y=>nx37624, A0=>label_5_output_8, A1=>nx42633, 
      A2=>nx41613);
   ix11643 : oai22 port map ( Y=>nx11642, A0=>nx37628, A1=>nx37641, B0=>
      max_calc_comparator_third_inp2_7, B1=>nx37636);
   ix26352 : oai21 port map ( Y=>nx26351, A0=>nx37632, A1=>nx41613, B0=>
      nx37634);
   max_calc_reg_comparator_third_inp2_7 : dff port map ( Q=>
      max_calc_comparator_third_inp2_7, QB=>nx37632, D=>nx26351, CLK=>clk);
   max_calc_reg_comparator_third_inp1_7 : dff port map ( Q=>
      max_calc_comparator_third_inp1_7, QB=>nx37636, D=>nx26361, CLK=>clk);
   ix26362 : oai21 port map ( Y=>nx26361, A0=>nx37636, A1=>nx41613, B0=>
      nx37639);
   ix37642 : aoi22 port map ( Y=>nx37641, A0=>nx37643, A1=>
      max_calc_comparator_third_inp1_6, B0=>nx11448, B1=>nx11626);
   max_calc_reg_comparator_third_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx37643, D=>nx26371, CLK=>clk);
   ix26372 : oai21 port map ( Y=>nx26371, A0=>nx37643, A1=>nx41613, B0=>
      nx37646);
   ix37647 : nand03 port map ( Y=>nx37646, A0=>label_6_output_6, A1=>nx42635, 
      A2=>nx41615);
   ix26382 : oai21 port map ( Y=>nx26381, A0=>nx37650, A1=>nx41615, B0=>
      nx37652);
   max_calc_reg_comparator_third_inp1_6 : dff port map ( Q=>
      max_calc_comparator_third_inp1_6, QB=>nx37650, D=>nx26381, CLK=>clk);
   ix37653 : nand03 port map ( Y=>nx37652, A0=>label_5_output_6, A1=>nx42635, 
      A2=>nx41615);
   ix11627 : oai22 port map ( Y=>nx11626, A0=>nx37656, A1=>nx37669, B0=>
      max_calc_comparator_third_inp2_5, B1=>nx37664);
   ix26392 : oai21 port map ( Y=>nx26391, A0=>nx37660, A1=>nx41615, B0=>
      nx37662);
   max_calc_reg_comparator_third_inp2_5 : dff port map ( Q=>
      max_calc_comparator_third_inp2_5, QB=>nx37660, D=>nx26391, CLK=>clk);
   max_calc_reg_comparator_third_inp1_5 : dff port map ( Q=>
      max_calc_comparator_third_inp1_5, QB=>nx37664, D=>nx26401, CLK=>clk);
   ix26402 : oai21 port map ( Y=>nx26401, A0=>nx37664, A1=>nx41615, B0=>
      nx37667);
   ix37670 : aoi22 port map ( Y=>nx37669, A0=>nx37671, A1=>
      max_calc_comparator_third_inp1_4, B0=>nx11492, B1=>nx11610);
   max_calc_reg_comparator_third_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx37671, D=>nx26411, CLK=>clk);
   ix26412 : oai21 port map ( Y=>nx26411, A0=>nx37671, A1=>nx41617, B0=>
      nx37674);
   ix37675 : nand03 port map ( Y=>nx37674, A0=>label_6_output_4, A1=>nx42635, 
      A2=>nx41617);
   ix26422 : oai21 port map ( Y=>nx26421, A0=>nx37678, A1=>nx41617, B0=>
      nx37680);
   max_calc_reg_comparator_third_inp1_4 : dff port map ( Q=>
      max_calc_comparator_third_inp1_4, QB=>nx37678, D=>nx26421, CLK=>clk);
   ix37681 : nand03 port map ( Y=>nx37680, A0=>label_5_output_4, A1=>nx42637, 
      A2=>nx41617);
   ix11611 : oai22 port map ( Y=>nx11610, A0=>nx37684, A1=>nx37697, B0=>
      max_calc_comparator_third_inp2_3, B1=>nx37692);
   ix26432 : oai21 port map ( Y=>nx26431, A0=>nx37688, A1=>nx41617, B0=>
      nx37690);
   max_calc_reg_comparator_third_inp2_3 : dff port map ( Q=>
      max_calc_comparator_third_inp2_3, QB=>nx37688, D=>nx26431, CLK=>clk);
   max_calc_reg_comparator_third_inp1_3 : dff port map ( Q=>
      max_calc_comparator_third_inp1_3, QB=>nx37692, D=>nx26441, CLK=>clk);
   ix26442 : oai21 port map ( Y=>nx26441, A0=>nx37692, A1=>nx41617, B0=>
      nx37695);
   ix37698 : aoi22 port map ( Y=>nx37697, A0=>nx37699, A1=>
      max_calc_comparator_third_inp1_2, B0=>nx11536, B1=>nx11594);
   max_calc_reg_comparator_third_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx37699, D=>nx26451, CLK=>clk);
   ix26452 : oai21 port map ( Y=>nx26451, A0=>nx37699, A1=>nx41619, B0=>
      nx37702);
   ix37703 : nand03 port map ( Y=>nx37702, A0=>label_6_output_2, A1=>nx42637, 
      A2=>nx41619);
   ix26462 : oai21 port map ( Y=>nx26461, A0=>nx37706, A1=>nx41619, B0=>
      nx37708);
   max_calc_reg_comparator_third_inp1_2 : dff port map ( Q=>
      max_calc_comparator_third_inp1_2, QB=>nx37706, D=>nx26461, CLK=>clk);
   ix37709 : nand03 port map ( Y=>nx37708, A0=>label_5_output_2, A1=>nx42637, 
      A2=>nx41619);
   ix11595 : oai21 port map ( Y=>nx11594, A0=>
      max_calc_comparator_third_inp2_1, A1=>nx37718, B0=>nx37723);
   ix26472 : oai21 port map ( Y=>nx26471, A0=>nx37714, A1=>nx41619, B0=>
      nx37716);
   max_calc_reg_comparator_third_inp2_1 : dff port map ( Q=>
      max_calc_comparator_third_inp2_1, QB=>nx37714, D=>nx26471, CLK=>clk);
   max_calc_reg_comparator_third_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx37718, D=>nx26481, CLK=>clk);
   ix26482 : oai21 port map ( Y=>nx26481, A0=>nx37718, A1=>nx41621, B0=>
      nx37721);
   ix37724 : oai21 port map ( Y=>nx37723, A0=>nx37725, A1=>
      max_calc_comparator_third_inp1_0, B0=>nx11558);
   max_calc_reg_comparator_third_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx37725, D=>nx26491, CLK=>clk);
   ix26492 : oai21 port map ( Y=>nx26491, A0=>nx37725, A1=>nx41621, B0=>
      nx37728);
   ix37729 : nand03 port map ( Y=>nx37728, A0=>label_6_output_0, A1=>nx42639, 
      A2=>nx41621);
   ix26502 : oai21 port map ( Y=>nx26501, A0=>nx37732, A1=>nx41621, B0=>
      nx37734);
   max_calc_reg_comparator_third_inp1_0 : dff port map ( Q=>
      max_calc_comparator_third_inp1_0, QB=>nx37732, D=>nx26501, CLK=>clk);
   ix37735 : nand03 port map ( Y=>nx37734, A0=>label_5_output_0, A1=>nx42639, 
      A2=>nx41621);
   ix26532 : oai21 port map ( Y=>nx26531, A0=>nx37740, A1=>nx41621, B0=>
      nx37742);
   max_calc_reg_comparator_third_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx37740, D=>nx26531, CLK=>clk);
   lat_label_6_input_15 : latch port map ( Q=>label_6_input_15, D=>nx11720, 
      CLK=>nx41691);
   reg_label_6_input_state_machine_15 : dffr port map ( Q=>
      label_6_input_state_machine_15, QB=>OPEN, D=>nx26511, CLK=>clk, R=>rst
   );
   ix11717 : xnor2 port map ( Y=>nx11716, A0=>nx37752, A1=>nx11714);
   ix37753 : aoi22 port map ( Y=>nx37752, A0=>label_6_output_14, A1=>
      booth_booth_integration_output_5_26, B0=>nx11242, B1=>nx11244);
   labelsregfile_label6_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_6_output_15, QB=>nx37756, D=>nx26521, CLK=>clk, R=>rst);
   ix26562 : oai21 port map ( Y=>nx26561, A0=>nx37760, A1=>nx41623, B0=>
      nx37762);
   max_calc_reg_comparator_third_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx37760, D=>nx26561, CLK=>clk);
   lat_label_5_input_15 : latch port map ( Q=>label_5_input_15, D=>nx11762, 
      CLK=>nx41691);
   reg_label_5_input_state_machine_15 : dffr port map ( Q=>
      label_5_input_state_machine_15, QB=>OPEN, D=>nx26541, CLK=>clk, R=>rst
   );
   ix11759 : xnor2 port map ( Y=>nx11758, A0=>nx37772, A1=>nx11756);
   ix37773 : aoi22 port map ( Y=>nx37772, A0=>label_5_output_14, A1=>
      booth_booth_integration_output_4_26, B0=>nx9924, B1=>nx9926);
   labelsregfile_label5_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_5_output_15, QB=>nx37776, D=>nx26551, CLK=>clk, R=>rst);
   ix29452 : oai21 port map ( Y=>nx29451, A0=>nx37785, A1=>nx41623, B0=>
      nx37787);
   max_calc_reg_comparator_second_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx37785, D=>nx29451, CLK=>clk);
   ix37788 : nand03 port map ( Y=>nx37787, A0=>nx42819, A1=>nx16298, A2=>
      nx41641);
   labelsregfile_label4_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_4_output_14, QB=>OPEN, D=>nx27411, CLK=>clk, R=>rst);
   lat_label_4_input_14 : latch port map ( Q=>label_4_input_14, D=>nx13114, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_14 : dffr port map ( Q=>
      label_4_input_state_machine_14, QB=>OPEN, D=>nx26591, CLK=>clk, R=>rst
   );
   ix13111 : xnor2 port map ( Y=>nx13110, A0=>nx13106, A1=>nx38415);
   ix13107 : oai22 port map ( Y=>nx13106, A0=>nx37799, A1=>nx38404, B0=>
      nx38414, B1=>nx38173);
   ix37800 : aoi22 port map ( Y=>nx37799, A0=>label_4_output_12, A1=>
      booth_booth_integration_output_3_24, B0=>nx13042, B1=>nx18499);
   labelsregfile_label4_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_4_output_12, QB=>OPEN, D=>nx27381, CLK=>clk, R=>rst);
   lat_label_4_input_12 : latch port map ( Q=>label_4_input_12, D=>nx13056, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_12 : dffr port map ( Q=>
      label_4_input_state_machine_12, QB=>OPEN, D=>nx27371, CLK=>clk, R=>rst
   );
   ix13053 : xnor2 port map ( Y=>nx13052, A0=>nx13042, A1=>nx38400);
   ix13043 : oai22 port map ( Y=>nx13042, A0=>nx37810, A1=>nx38389, B0=>
      nx38399, B1=>nx38137);
   ix37811 : aoi22 port map ( Y=>nx37810, A0=>label_4_output_10, A1=>
      booth_booth_integration_output_3_22, B0=>nx12978, B1=>nx18497);
   labelsregfile_label4_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_4_output_10, QB=>OPEN, D=>nx27341, CLK=>clk, R=>rst);
   lat_label_4_input_10 : latch port map ( Q=>label_4_input_10, D=>nx12992, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_10 : dffr port map ( Q=>
      label_4_input_state_machine_10, QB=>OPEN, D=>nx27331, CLK=>clk, R=>rst
   );
   ix12989 : xnor2 port map ( Y=>nx12988, A0=>nx12978, A1=>nx38385);
   ix12979 : oai22 port map ( Y=>nx12978, A0=>nx37821, A1=>nx38374, B0=>
      nx38384, B1=>nx38101);
   ix37822 : aoi22 port map ( Y=>nx37821, A0=>label_4_output_8, A1=>
      booth_booth_integration_output_3_20, B0=>nx12914, B1=>nx18493);
   labelsregfile_label4_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_4_output_8, QB=>OPEN, D=>nx27301, CLK=>clk, R=>rst);
   lat_label_4_input_8 : latch port map ( Q=>label_4_input_8, D=>nx12928, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_8 : dffr port map ( Q=>
      label_4_input_state_machine_8, QB=>OPEN, D=>nx27291, CLK=>clk, R=>rst
   );
   ix12925 : xnor2 port map ( Y=>nx12924, A0=>nx12914, A1=>nx38370);
   ix12915 : oai22 port map ( Y=>nx12914, A0=>nx37832, A1=>nx38359, B0=>
      nx38369, B1=>nx38063);
   ix37833 : aoi22 port map ( Y=>nx37832, A0=>label_4_output_6, A1=>
      booth_booth_integration_output_3_18, B0=>nx12850, B1=>nx18490);
   labelsregfile_label4_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_4_output_6, QB=>OPEN, D=>nx27261, CLK=>clk, R=>rst);
   lat_label_4_input_6 : latch port map ( Q=>label_4_input_6, D=>nx12864, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_6 : dffr port map ( Q=>
      label_4_input_state_machine_6, QB=>OPEN, D=>nx27251, CLK=>clk, R=>rst
   );
   ix12861 : xnor2 port map ( Y=>nx12860, A0=>nx12850, A1=>nx38355);
   ix12851 : oai22 port map ( Y=>nx12850, A0=>nx37843, A1=>nx38344, B0=>
      nx38354, B1=>nx38024);
   ix37844 : aoi22 port map ( Y=>nx37843, A0=>label_4_output_4, A1=>
      booth_booth_integration_output_3_16, B0=>nx12786, B1=>nx18488);
   labelsregfile_label4_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_4_output_4, QB=>OPEN, D=>nx27221, CLK=>clk, R=>rst);
   lat_label_4_input_4 : latch port map ( Q=>label_4_input_4, D=>nx12800, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_4 : dffr port map ( Q=>
      label_4_input_state_machine_4, QB=>OPEN, D=>nx27211, CLK=>clk, R=>rst
   );
   ix12797 : xnor2 port map ( Y=>nx12796, A0=>nx12786, A1=>nx38340);
   ix12787 : oai22 port map ( Y=>nx12786, A0=>nx37854, A1=>nx38329, B0=>
      nx38339, B1=>nx38307);
   ix37855 : aoi22 port map ( Y=>nx37854, A0=>label_4_output_2, A1=>
      booth_booth_integration_output_3_14, B0=>nx12722, B1=>nx18486);
   labelsregfile_label4_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_4_output_2, QB=>OPEN, D=>nx27181, CLK=>clk, R=>rst);
   lat_label_4_input_2 : latch port map ( Q=>label_4_input_2, D=>nx12736, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_2 : dffr port map ( Q=>
      label_4_input_state_machine_2, QB=>OPEN, D=>nx27171, CLK=>clk, R=>rst
   );
   ix12733 : xnor2 port map ( Y=>nx12732, A0=>nx12722, A1=>nx38325);
   ix12723 : oai22 port map ( Y=>nx12722, A0=>nx37865, A1=>nx38314, B0=>
      nx38324, B1=>nx38310);
   ix37866 : nand02 port map ( Y=>nx37865, A0=>label_4_output_0, A1=>
      booth_booth_integration_output_3_12);
   labelsregfile_label4_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_4_output_0, QB=>OPEN, D=>nx27141, CLK=>clk, R=>rst);
   lat_label_4_input_0 : latch port map ( Q=>label_4_input_0, D=>nx12678, 
      CLK=>nx41691);
   ix12679 : oai21 port map ( Y=>nx12678, A0=>nx37871, A1=>nx41453, B0=>
      nx37875);
   reg_label_4_input_state_machine_0 : dffr port map ( Q=>
      label_4_input_state_machine_0, QB=>nx37871, D=>nx27131, CLK=>clk, R=>
      rst);
   ix37876 : oai21 port map ( Y=>nx37875, A0=>
      booth_booth_integration_output_3_12, A1=>label_4_output_0, B0=>nx12666
   );
   booth_booth_integrtaion_3_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_12, QB=>OPEN, D=>nx27121, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_13, QB=>nx38310, D=>nx27111, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_14, QB=>OPEN, D=>nx27101, CLK=>clk, R
      =>rst);
   ix37889 : aoi22 port map ( Y=>nx37888, A0=>nx41797, A1=>nx42055, B0=>
      nx12608, B1=>nx12614);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_reg_output_0, QB=>OPEN, 
      D=>nx26621, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_0, QB=>OPEN, D=>nx26607, CLK
      =>clk, S=>nx41499);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_reg_output_9, QB=>OPEN, 
      D=>nx26801, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_9, QB=>OPEN, D=>nx26791, CLK
      =>clk, R=>nx41499);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12772, QB=>OPEN, D=>nx26781, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_8, QB=>OPEN, D=>nx26771, CLK
      =>clk, R=>nx41499);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12773, QB=>OPEN, D=>nx26761, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_7, QB=>OPEN, D=>nx26751, CLK
      =>clk, R=>nx41499);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12774, QB=>OPEN, D=>nx26741, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_6, QB=>OPEN, D=>nx26731, CLK
      =>clk, R=>nx41497);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12775, QB=>OPEN, D=>nx26721, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_5, QB=>OPEN, D=>nx26711, CLK
      =>clk, R=>nx41497);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12776, QB=>OPEN, D=>nx26701, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_4, QB=>OPEN, D=>nx26691, CLK
      =>clk, R=>nx41497);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12777, QB=>OPEN, D=>nx26681, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_3, QB=>OPEN, D=>nx26671, CLK
      =>clk, R=>nx41497);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12778, QB=>OPEN, D=>nx26661, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_2, QB=>OPEN, D=>nx26651, CLK
      =>clk, R=>nx41497);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12779, QB=>OPEN, D=>nx26641, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_1, QB=>OPEN, D=>nx26631, CLK
      =>clk, R=>nx41497);
   ix26602 : nand02 port map ( Y=>nx26601, A0=>nx42953, A1=>nx42041);
   booth_booth_integrtaion_3_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx37935, D=>nx26601, CLK=>clk, S=>nx41497);
   ix12609 : nand02 port map ( Y=>nx12608, A0=>nx37956, A1=>nx38014);
   ix37957 : oai21 port map ( Y=>nx37956, A0=>nx42067, A1=>nx42063, B0=>
      data_in(48));
   ix26932 : oai21 port map ( Y=>nx26931, A0=>nx37961, A1=>nx42697, B0=>
      nx37963);
   booth_booth_integrtaion_3_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx37961, D=>nx26931, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12168, QB=>nx38012, D=>nx26921, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12167, QB=>OPEN, D=>nx26911, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12166, QB=>OPEN, D=>nx26901, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12165, QB=>OPEN, D=>nx26891, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12164, QB=>OPEN, D=>nx26881, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12163, QB=>OPEN, D=>nx26871, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12162, QB=>OPEN, D=>nx26861, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12161, QB=>OPEN, D=>nx26851, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12160, QB=>OPEN, D=>nx26841, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12159, QB=>OPEN, D=>nx26831, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12158, QB=>OPEN, D=>nx26821, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12157, QB=>OPEN, D=>nx26811, CLK=>clk, R=>rst);
   ix38019 : xnor2 port map ( Y=>nx38018, A0=>nx12078, A1=>nx18461);
   ix27072 : oai21 port map ( Y=>nx27071, A0=>nx38024, A1=>nx42697, B0=>
      nx38026);
   booth_booth_integrtaion_3_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_17, QB=>nx38024, D=>nx27071, CLK=>clk, 
      R=>rst);
   ix38027 : nand03 port map ( Y=>nx38026, A0=>nx42705, A1=>nx12586, A2=>
      nx42701);
   ix12587 : xnor2 port map ( Y=>nx12586, A0=>nx38029, A1=>nx18463);
   ix38030 : aoi22 port map ( Y=>nx38029, A0=>
      booth_booth_integration_output_3_17, A1=>nx12102, B0=>nx12078, B1=>
      nx18461);
   ix12093 : nor02_2x port map ( Y=>nx12092, A0=>data_in(48), A1=>
      data_in(49));
   ix27062 : oai21 port map ( Y=>nx27061, A0=>nx38044, A1=>nx42697, B0=>
      nx38046);
   booth_booth_integrtaion_3_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_18, QB=>nx38044, D=>nx27061, CLK=>clk, 
      R=>rst);
   ix38047 : nand03 port map ( Y=>nx38046, A0=>nx42705, A1=>nx12574, A2=>
      nx42701);
   ix12575 : xnor2 port map ( Y=>nx12574, A0=>nx12130, A1=>nx38059);
   ix12131 : oai22 port map ( Y=>nx12130, A0=>nx38029, A1=>nx38050, B0=>
      nx38044, B1=>nx42709);
   ix38053 : aoi32 port map ( Y=>nx38052, A0=>nx12112, A1=>nx42067, A2=>
      nx38055, B0=>data_in(50), B1=>nx42063);
   ix12113 : oai21 port map ( Y=>nx12112, A0=>data_in(48), A1=>data_in(49), 
      B0=>data_in(50));
   ix27052 : oai21 port map ( Y=>nx27051, A0=>nx38063, A1=>nx42697, B0=>
      nx38065);
   booth_booth_integrtaion_3_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_19, QB=>nx38063, D=>nx27051, CLK=>clk, 
      R=>rst);
   ix38066 : nand03 port map ( Y=>nx38065, A0=>nx42705, A1=>nx12562, A2=>
      nx42701);
   ix12563 : xnor2 port map ( Y=>nx12562, A0=>nx38068, A1=>nx18467);
   ix38069 : aoi22 port map ( Y=>nx38068, A0=>
      booth_booth_integration_output_3_19, A1=>nx12150, B0=>nx12130, B1=>
      nx18465);
   ix12151 : oai32 port map ( Y=>nx12150, A0=>nx38071, A1=>nx38034, A2=>
      nx12140, B0=>nx38074, B1=>nx38039);
   ix12117 : nor03_2x port map ( Y=>nx12116, A0=>data_in(50), A1=>
      data_in(48), A2=>data_in(49));
   ix38075 : inv01 port map ( Y=>nx38074, A=>data_in(51));
   ix12141 : nor04 port map ( Y=>nx12140, A0=>data_in(51), A1=>data_in(50), 
      A2=>data_in(48), A3=>data_in(49));
   ix38083 : xnor2 port map ( Y=>nx38082, A0=>nx12178, A1=>nx18469);
   ix12179 : oai22 port map ( Y=>nx12178, A0=>nx38068, A1=>nx38085, B0=>
      nx38096, B1=>nx42711);
   ix38088 : aoi32 port map ( Y=>nx38087, A0=>nx12160, A1=>nx42067, A2=>
      nx38092, B0=>data_in(52), B1=>nx42063);
   ix12161 : nand02 port map ( Y=>nx12160, A0=>nx38090, A1=>data_in(52));
   ix38093 : nand02 port map ( Y=>nx38092, A0=>nx38094, A1=>nx12140);
   ix38095 : inv01 port map ( Y=>nx38094, A=>data_in(52));
   booth_booth_integrtaion_3_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_20, QB=>nx38096, D=>nx27041, CLK=>clk, 
      R=>rst);
   ix27032 : oai21 port map ( Y=>nx27031, A0=>nx38101, A1=>nx42697, B0=>
      nx38103);
   booth_booth_integrtaion_3_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_21, QB=>nx38101, D=>nx27031, CLK=>clk, 
      R=>rst);
   ix38104 : nand03 port map ( Y=>nx38103, A0=>nx42705, A1=>nx12538, A2=>
      nx42701);
   ix12539 : xnor2 port map ( Y=>nx12538, A0=>nx38106, A1=>nx18471);
   ix38107 : aoi22 port map ( Y=>nx38106, A0=>
      booth_booth_integration_output_3_21, A1=>nx12198, B0=>nx12178, B1=>
      nx18469);
   ix12189 : nor02_2x port map ( Y=>nx12188, A0=>data_in(53), A1=>nx38092);
   ix38119 : xnor2 port map ( Y=>nx38118, A0=>nx12226, A1=>nx18472);
   ix12227 : oai22 port map ( Y=>nx12226, A0=>nx38106, A1=>nx38121, B0=>
      nx38132, B1=>nx42713);
   ix38124 : aoi32 port map ( Y=>nx38123, A0=>nx12208, A1=>nx42067, A2=>
      nx38128, B0=>data_in(54), B1=>nx42063);
   ix12209 : nand02 port map ( Y=>nx12208, A0=>nx38126, A1=>data_in(54));
   ix38129 : nand02 port map ( Y=>nx38128, A0=>nx38130, A1=>nx12188);
   ix38131 : inv01 port map ( Y=>nx38130, A=>data_in(54));
   booth_booth_integrtaion_3_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_22, QB=>nx38132, D=>nx27021, CLK=>clk, 
      R=>rst);
   ix27012 : oai21 port map ( Y=>nx27011, A0=>nx38137, A1=>nx42699, B0=>
      nx38139);
   booth_booth_integrtaion_3_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_23, QB=>nx38137, D=>nx27011, CLK=>clk, 
      R=>rst);
   ix38140 : nand03 port map ( Y=>nx38139, A0=>nx42705, A1=>nx12514, A2=>
      nx42701);
   ix12515 : xnor2 port map ( Y=>nx12514, A0=>nx38142, A1=>nx18473);
   ix38143 : aoi22 port map ( Y=>nx38142, A0=>
      booth_booth_integration_output_3_23, A1=>nx12246, B0=>nx12226, B1=>
      nx18472);
   ix12237 : nor02_2x port map ( Y=>nx12236, A0=>data_in(55), A1=>nx38128);
   ix38155 : xnor2 port map ( Y=>nx38154, A0=>nx12274, A1=>nx18474);
   ix12275 : oai22 port map ( Y=>nx12274, A0=>nx38142, A1=>nx38157, B0=>
      nx38168, B1=>nx42715);
   ix38160 : aoi32 port map ( Y=>nx38159, A0=>nx12256, A1=>nx42067, A2=>
      nx38164, B0=>data_in(56), B1=>nx42063);
   ix12257 : nand02 port map ( Y=>nx12256, A0=>nx38162, A1=>data_in(56));
   ix38165 : nand02 port map ( Y=>nx38164, A0=>nx38166, A1=>nx12236);
   ix38167 : inv01 port map ( Y=>nx38166, A=>data_in(56));
   booth_booth_integrtaion_3_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_24, QB=>nx38168, D=>nx27001, CLK=>clk, 
      R=>rst);
   ix26992 : oai21 port map ( Y=>nx26991, A0=>nx38173, A1=>nx42699, B0=>
      nx38175);
   booth_booth_integrtaion_3_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_25, QB=>nx38173, D=>nx26991, CLK=>clk, 
      R=>rst);
   ix38176 : nand03 port map ( Y=>nx38175, A0=>nx42705, A1=>nx12490, A2=>
      nx42701);
   ix12491 : xnor2 port map ( Y=>nx12490, A0=>nx38178, A1=>nx18475);
   ix38179 : aoi22 port map ( Y=>nx38178, A0=>
      booth_booth_integration_output_3_25, A1=>nx12294, B0=>nx12274, B1=>
      nx18474);
   ix12285 : nor02_2x port map ( Y=>nx12284, A0=>data_in(57), A1=>nx38164);
   ix38191 : xnor2 port map ( Y=>nx38190, A0=>nx12322, A1=>nx18476);
   ix12323 : oai22 port map ( Y=>nx12322, A0=>nx38178, A1=>nx38193, B0=>
      nx38204, B1=>nx42717);
   ix38196 : aoi32 port map ( Y=>nx38195, A0=>nx12304, A1=>nx42067, A2=>
      nx38200, B0=>data_in(58), B1=>nx42063);
   ix12305 : nand02 port map ( Y=>nx12304, A0=>nx38198, A1=>data_in(58));
   ix38201 : nand02 port map ( Y=>nx38200, A0=>nx38202, A1=>nx12284);
   ix38203 : inv01 port map ( Y=>nx38202, A=>data_in(58));
   booth_booth_integrtaion_3_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_26, QB=>nx38204, D=>nx26981, CLK=>clk, 
      R=>rst);
   ix26972 : oai21 port map ( Y=>nx26971, A0=>nx38209, A1=>nx42699, B0=>
      nx38211);
   booth_booth_integrtaion_3_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_27, QB=>nx38209, D=>nx26971, CLK=>clk, 
      R=>rst);
   ix38212 : nand03 port map ( Y=>nx38211, A0=>nx43299, A1=>nx12466, A2=>
      nx42701);
   ix12467 : xnor2 port map ( Y=>nx12466, A0=>nx38214, A1=>nx18477);
   ix38215 : aoi22 port map ( Y=>nx38214, A0=>
      booth_booth_integration_output_3_27, A1=>nx12342, B0=>nx12322, B1=>
      nx18476);
   ix12333 : nor02_2x port map ( Y=>nx12332, A0=>data_in(59), A1=>nx38200);
   ix38227 : xnor2 port map ( Y=>nx38226, A0=>nx12370, A1=>nx18479);
   ix12371 : oai22 port map ( Y=>nx12370, A0=>nx38214, A1=>nx38229, B0=>
      nx38240, B1=>nx42719);
   ix38232 : aoi32 port map ( Y=>nx38231, A0=>nx12352, A1=>nx42069, A2=>
      nx38236, B0=>data_in(60), B1=>nx42063);
   ix12353 : nand02 port map ( Y=>nx12352, A0=>nx38234, A1=>data_in(60));
   ix38237 : nand02 port map ( Y=>nx38236, A0=>nx38238, A1=>nx12332);
   ix38239 : inv01 port map ( Y=>nx38238, A=>data_in(60));
   booth_booth_integrtaion_3_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12156, QB=>nx38240, D=>nx26961, CLK=>clk, R=>rst);
   ix26952 : oai21 port map ( Y=>nx26951, A0=>nx38245, A1=>nx42699, B0=>
      nx38247);
   booth_booth_integrtaion_3_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12155, QB=>nx38245, D=>nx26951, CLK=>clk, R=>rst);
   ix38248 : nand03 port map ( Y=>nx38247, A0=>nx43299, A1=>nx12442, A2=>
      nx42699);
   ix12443 : xnor2 port map ( Y=>nx12442, A0=>nx38250, A1=>nx18481);
   ix38251 : aoi22 port map ( Y=>nx38250, A0=>booth_output_29_dup_12155, A1
      =>nx12390, B0=>nx12370, B1=>nx18479);
   ix12381 : nor02_2x port map ( Y=>nx12380, A0=>data_in(61), A1=>nx38236);
   ix26942 : oai21 port map ( Y=>nx26941, A0=>nx38261, A1=>nx42699, B0=>
      nx38263);
   booth_booth_integrtaion_3_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx38261, D=>nx26941, CLK=>clk, R=>rst);
   ix38264 : nand03 port map ( Y=>nx38263, A0=>nx43299, A1=>nx12430, A2=>
      nx42699);
   ix12431 : xnor2 port map ( Y=>nx12430, A0=>nx12418, A1=>nx38278);
   ix12419 : oai22 port map ( Y=>nx12418, A0=>nx38250, A1=>nx38267, B0=>
      nx38261, B1=>nx42721);
   ix38270 : aoi32 port map ( Y=>nx38269, A0=>nx12400, A1=>nx42069, A2=>
      nx38274, B0=>data_in(62), B1=>nx42065);
   ix12401 : nand02 port map ( Y=>nx12400, A0=>nx38272, A1=>data_in(62));
   ix38275 : nand02 port map ( Y=>nx38274, A0=>nx38276, A1=>nx12380);
   ix38277 : inv01 port map ( Y=>nx38276, A=>data_in(62));
   ix12427 : oai22 port map ( Y=>nx12426, A0=>nx38034, A1=>nx38281, B0=>
      nx38283, B1=>nx38039);
   ix38282 : xnor2 port map ( Y=>nx38281, A0=>data_in(63), A1=>nx38274);
   ix38284 : inv01 port map ( Y=>nx38283, A=>data_in(63));
   ix38286 : aoi32 port map ( Y=>nx38285, A0=>nx12376, A1=>nx42069, A2=>
      nx38272, B0=>data_in(61), B1=>nx42065);
   ix12377 : nand02 port map ( Y=>nx12376, A0=>nx38236, A1=>data_in(61));
   ix38289 : aoi32 port map ( Y=>nx38288, A0=>nx12328, A1=>nx42069, A2=>
      nx38234, B0=>data_in(59), B1=>nx42065);
   ix12329 : nand02 port map ( Y=>nx12328, A0=>nx38200, A1=>data_in(59));
   ix38292 : aoi32 port map ( Y=>nx38291, A0=>nx12280, A1=>nx42069, A2=>
      nx38198, B0=>data_in(57), B1=>nx42065);
   ix12281 : nand02 port map ( Y=>nx12280, A0=>nx38164, A1=>data_in(57));
   ix38295 : aoi32 port map ( Y=>nx38294, A0=>nx12232, A1=>nx42069, A2=>
      nx38162, B0=>data_in(55), B1=>nx42065);
   ix12233 : nand02 port map ( Y=>nx12232, A0=>nx38128, A1=>data_in(55));
   ix38298 : aoi32 port map ( Y=>nx38297, A0=>nx12184, A1=>nx42071, A2=>
      nx38126, B0=>data_in(53), B1=>nx42065);
   ix12185 : nand02 port map ( Y=>nx12184, A0=>nx38092, A1=>data_in(53));
   ix38301 : aoi32 port map ( Y=>nx38300, A0=>nx12086, A1=>nx42071, A2=>
      nx38303, B0=>data_in(49), B1=>nx42065);
   ix12087 : nand02 port map ( Y=>nx12086, A0=>data_in(49), A1=>data_in(48)
   );
   booth_booth_integrtaion_3_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_16, QB=>nx38014, D=>nx27081, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_15, QB=>nx38307, D=>nx27091, CLK=>clk, 
      R=>rst);
   ix12667 : aoi21 port map ( Y=>nx12666, A0=>label_4_output_0, A1=>
      booth_booth_integration_output_3_12, B0=>nx43055);
   labelsregfile_label4_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_4_output_1, QB=>nx38324, D=>nx27161, CLK=>clk, R=>rst);
   lat_label_4_input_1 : latch port map ( Q=>label_4_input_1, D=>nx12704, 
      CLK=>nx41691);
   reg_label_4_input_state_machine_1 : dffr port map ( Q=>
      label_4_input_state_machine_1, QB=>OPEN, D=>nx27151, CLK=>clk, R=>rst
   );
   ix12701 : xor2 port map ( Y=>nx12700, A0=>nx37865, A1=>nx38314);
   ix38326 : xnor2 port map ( Y=>nx38325, A0=>
      booth_booth_integration_output_3_14, A1=>label_4_output_2);
   labelsregfile_label4_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_4_output_3, QB=>nx38339, D=>nx27201, CLK=>clk, R=>rst);
   lat_label_4_input_3 : latch port map ( Q=>label_4_input_3, D=>nx12768, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_3 : dffr port map ( Q=>
      label_4_input_state_machine_3, QB=>OPEN, D=>nx27191, CLK=>clk, R=>rst
   );
   ix12765 : xor2 port map ( Y=>nx12764, A0=>nx37854, A1=>nx38329);
   labelsregfile_label4_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_4_output_5, QB=>nx38354, D=>nx27241, CLK=>clk, R=>rst);
   lat_label_4_input_5 : latch port map ( Q=>label_4_input_5, D=>nx12832, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_5 : dffr port map ( Q=>
      label_4_input_state_machine_5, QB=>OPEN, D=>nx27231, CLK=>clk, R=>rst
   );
   ix12829 : xor2 port map ( Y=>nx12828, A0=>nx37843, A1=>nx38344);
   labelsregfile_label4_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_4_output_7, QB=>nx38369, D=>nx27281, CLK=>clk, R=>rst);
   lat_label_4_input_7 : latch port map ( Q=>label_4_input_7, D=>nx12896, 
      CLK=>nx41693);
   reg_label_4_input_state_machine_7 : dffr port map ( Q=>
      label_4_input_state_machine_7, QB=>OPEN, D=>nx27271, CLK=>clk, R=>rst
   );
   ix12893 : xor2 port map ( Y=>nx12892, A0=>nx37832, A1=>nx38359);
   labelsregfile_label4_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_4_output_9, QB=>nx38384, D=>nx27321, CLK=>clk, R=>rst);
   lat_label_4_input_9 : latch port map ( Q=>label_4_input_9, D=>nx12960, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_9 : dffr port map ( Q=>
      label_4_input_state_machine_9, QB=>OPEN, D=>nx27311, CLK=>clk, R=>rst
   );
   ix12957 : xor2 port map ( Y=>nx12956, A0=>nx37821, A1=>nx38374);
   labelsregfile_label4_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_4_output_11, QB=>nx38399, D=>nx27361, CLK=>clk, R=>rst);
   lat_label_4_input_11 : latch port map ( Q=>label_4_input_11, D=>nx13024, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_11 : dffr port map ( Q=>
      label_4_input_state_machine_11, QB=>OPEN, D=>nx27351, CLK=>clk, R=>rst
   );
   ix13021 : xor2 port map ( Y=>nx13020, A0=>nx37810, A1=>nx38389);
   labelsregfile_label4_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_4_output_13, QB=>nx38414, D=>nx27401, CLK=>clk, R=>rst);
   lat_label_4_input_13 : latch port map ( Q=>label_4_input_13, D=>nx13088, 
      CLK=>nx41695);
   reg_label_4_input_state_machine_13 : dffr port map ( Q=>
      label_4_input_state_machine_13, QB=>OPEN, D=>nx27391, CLK=>clk, R=>rst
   );
   ix13085 : xor2 port map ( Y=>nx13084, A0=>nx37799, A1=>nx38404);
   max_calc_reg_ans4_14 : dff port map ( Q=>max_calc_ans4_14, QB=>OPEN, D=>
      nx29441, CLK=>clk);
   ix29442 : ao32 port map ( Y=>nx29441, A0=>nx42819, A1=>nx16284, A2=>
      nx41811, B0=>max_calc_ans4_14, B1=>nx42679);
   ix28252 : oai21 port map ( Y=>nx28251, A0=>nx38423, A1=>nx41623, B0=>
      nx38425);
   max_calc_reg_comparator_fourth_inp1_14 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_14, QB=>nx38423, D=>nx28251, CLK=>clk
   );
   ix38426 : nand03 port map ( Y=>nx38425, A0=>label_7_output_14, A1=>
      nx42639, A2=>nx41623);
   labelsregfile_label7_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_7_output_14, QB=>OPEN, D=>nx28241, CLK=>clk, R=>rst);
   lat_label_7_input_14 : latch port map ( Q=>label_7_input_14, D=>nx14424, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_14 : dffr port map ( Q=>
      label_7_input_state_machine_14, QB=>OPEN, D=>nx27421, CLK=>clk, R=>rst
   );
   ix14421 : xnor2 port map ( Y=>nx14420, A0=>nx14416, A1=>nx39052);
   ix14417 : oai22 port map ( Y=>nx14416, A0=>nx38436, A1=>nx39041, B0=>
      nx39051, B1=>nx38810);
   ix38437 : aoi22 port map ( Y=>nx38436, A0=>label_7_output_12, A1=>
      booth_booth_integration_output_6_24, B0=>nx14352, B1=>nx18539);
   labelsregfile_label7_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_7_output_12, QB=>OPEN, D=>nx28211, CLK=>clk, R=>rst);
   lat_label_7_input_12 : latch port map ( Q=>label_7_input_12, D=>nx14366, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_12 : dffr port map ( Q=>
      label_7_input_state_machine_12, QB=>OPEN, D=>nx28201, CLK=>clk, R=>rst
   );
   ix14363 : xnor2 port map ( Y=>nx14362, A0=>nx14352, A1=>nx39037);
   ix14353 : oai22 port map ( Y=>nx14352, A0=>nx38447, A1=>nx39026, B0=>
      nx39036, B1=>nx38774);
   ix38448 : aoi22 port map ( Y=>nx38447, A0=>label_7_output_10, A1=>
      booth_booth_integration_output_6_22, B0=>nx14288, B1=>nx18535);
   labelsregfile_label7_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_7_output_10, QB=>OPEN, D=>nx28171, CLK=>clk, R=>rst);
   lat_label_7_input_10 : latch port map ( Q=>label_7_input_10, D=>nx14302, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_10 : dffr port map ( Q=>
      label_7_input_state_machine_10, QB=>OPEN, D=>nx28161, CLK=>clk, R=>rst
   );
   ix14299 : xnor2 port map ( Y=>nx14298, A0=>nx14288, A1=>nx39022);
   ix14289 : oai22 port map ( Y=>nx14288, A0=>nx38458, A1=>nx39011, B0=>
      nx39021, B1=>nx38738);
   ix38459 : aoi22 port map ( Y=>nx38458, A0=>label_7_output_8, A1=>
      booth_booth_integration_output_6_20, B0=>nx14224, B1=>nx18531);
   labelsregfile_label7_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_7_output_8, QB=>OPEN, D=>nx28131, CLK=>clk, R=>rst);
   lat_label_7_input_8 : latch port map ( Q=>label_7_input_8, D=>nx14238, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_8 : dffr port map ( Q=>
      label_7_input_state_machine_8, QB=>OPEN, D=>nx28121, CLK=>clk, R=>rst
   );
   ix14235 : xnor2 port map ( Y=>nx14234, A0=>nx14224, A1=>nx39007);
   ix14225 : oai22 port map ( Y=>nx14224, A0=>nx38469, A1=>nx38996, B0=>
      nx39006, B1=>nx38700);
   ix38470 : aoi22 port map ( Y=>nx38469, A0=>label_7_output_6, A1=>
      booth_booth_integration_output_6_18, B0=>nx14160, B1=>nx18528);
   labelsregfile_label7_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_7_output_6, QB=>OPEN, D=>nx28091, CLK=>clk, R=>rst);
   lat_label_7_input_6 : latch port map ( Q=>label_7_input_6, D=>nx14174, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_6 : dffr port map ( Q=>
      label_7_input_state_machine_6, QB=>OPEN, D=>nx28081, CLK=>clk, R=>rst
   );
   ix14171 : xnor2 port map ( Y=>nx14170, A0=>nx14160, A1=>nx38992);
   ix14161 : oai22 port map ( Y=>nx14160, A0=>nx38480, A1=>nx38981, B0=>
      nx38991, B1=>nx38661);
   ix38481 : aoi22 port map ( Y=>nx38480, A0=>label_7_output_4, A1=>
      booth_booth_integration_output_6_16, B0=>nx14096, B1=>nx18526);
   labelsregfile_label7_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_7_output_4, QB=>OPEN, D=>nx28051, CLK=>clk, R=>rst);
   lat_label_7_input_4 : latch port map ( Q=>label_7_input_4, D=>nx14110, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_4 : dffr port map ( Q=>
      label_7_input_state_machine_4, QB=>OPEN, D=>nx28041, CLK=>clk, R=>rst
   );
   ix14107 : xnor2 port map ( Y=>nx14106, A0=>nx14096, A1=>nx38977);
   ix14097 : oai22 port map ( Y=>nx14096, A0=>nx38491, A1=>nx38966, B0=>
      nx38976, B1=>nx38944);
   ix38492 : aoi22 port map ( Y=>nx38491, A0=>label_7_output_2, A1=>
      booth_booth_integration_output_6_14, B0=>nx14032, B1=>nx18524);
   labelsregfile_label7_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_7_output_2, QB=>OPEN, D=>nx28011, CLK=>clk, R=>rst);
   lat_label_7_input_2 : latch port map ( Q=>label_7_input_2, D=>nx14046, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_2 : dffr port map ( Q=>
      label_7_input_state_machine_2, QB=>OPEN, D=>nx28001, CLK=>clk, R=>rst
   );
   ix14043 : xnor2 port map ( Y=>nx14042, A0=>nx14032, A1=>nx38962);
   ix14033 : oai22 port map ( Y=>nx14032, A0=>nx38502, A1=>nx38951, B0=>
      nx38961, B1=>nx38947);
   ix38503 : nand02 port map ( Y=>nx38502, A0=>label_7_output_0, A1=>
      booth_booth_integration_output_6_12);
   labelsregfile_label7_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_7_output_0, QB=>OPEN, D=>nx27971, CLK=>clk, R=>rst);
   lat_label_7_input_0 : latch port map ( Q=>label_7_input_0, D=>nx13988, 
      CLK=>nx41695);
   ix13989 : oai21 port map ( Y=>nx13988, A0=>nx38508, A1=>nx41457, B0=>
      nx38512);
   reg_label_7_input_state_machine_0 : dffr port map ( Q=>
      label_7_input_state_machine_0, QB=>nx38508, D=>nx27961, CLK=>clk, R=>
      rst);
   ix38513 : oai21 port map ( Y=>nx38512, A0=>
      booth_booth_integration_output_6_12, A1=>label_7_output_0, B0=>nx13976
   );
   booth_booth_integrtaion_6_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_12, QB=>OPEN, D=>nx27951, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_13, QB=>nx38947, D=>nx27941, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_14, QB=>OPEN, D=>nx27931, CLK=>clk, R
      =>rst);
   ix38526 : aoi22 port map ( Y=>nx38525, A0=>nx41797, A1=>nx42087, B0=>
      nx13918, B1=>nx13924);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_reg_output_0, QB=>OPEN, 
      D=>nx27451, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_0, QB=>OPEN, D=>nx27437, CLK
      =>clk, S=>nx41503);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_reg_output_9, QB=>OPEN, 
      D=>nx27631, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_9, QB=>OPEN, D=>nx27621, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12856, QB=>OPEN, D=>nx27611, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_8, QB=>OPEN, D=>nx27601, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12857, QB=>OPEN, D=>nx27591, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_7, QB=>OPEN, D=>nx27581, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12858, QB=>OPEN, D=>nx27571, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_6, QB=>OPEN, D=>nx27561, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12859, QB=>OPEN, D=>nx27551, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_5, QB=>OPEN, D=>nx27541, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12860, QB=>OPEN, D=>nx27531, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_4, QB=>OPEN, D=>nx27521, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12861, QB=>OPEN, D=>nx27511, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_3, QB=>OPEN, D=>nx27501, CLK
      =>clk, R=>nx41501);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12862, QB=>OPEN, D=>nx27491, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_2, QB=>OPEN, D=>nx27481, CLK
      =>clk, R=>nx41499);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12863, QB=>OPEN, D=>nx27471, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_1, QB=>OPEN, D=>nx27461, CLK
      =>clk, R=>nx41499);
   ix27432 : nand02 port map ( Y=>nx27431, A0=>nx42957, A1=>nx42073);
   booth_booth_integrtaion_6_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx38572, D=>nx27431, CLK=>clk, S=>nx41499);
   ix13919 : nand02 port map ( Y=>nx13918, A0=>nx38593, A1=>nx38651);
   ix38594 : oai21 port map ( Y=>nx38593, A0=>nx42099, A1=>nx42095, B0=>
      data_in(96));
   ix27762 : oai21 port map ( Y=>nx27761, A0=>nx38598, A1=>nx42723, B0=>
      nx38600);
   booth_booth_integrtaion_6_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx38598, D=>nx27761, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12225, QB=>nx38649, D=>nx27751, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12224, QB=>OPEN, D=>nx27741, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12223, QB=>OPEN, D=>nx27731, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12222, QB=>OPEN, D=>nx27721, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12221, QB=>OPEN, D=>nx27711, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12220, QB=>OPEN, D=>nx27701, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12219, QB=>OPEN, D=>nx27691, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12218, QB=>OPEN, D=>nx27681, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12217, QB=>OPEN, D=>nx27671, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12216, QB=>OPEN, D=>nx27661, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12215, QB=>OPEN, D=>nx27651, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12214, QB=>OPEN, D=>nx27641, CLK=>clk, R=>rst);
   ix38656 : xnor2 port map ( Y=>nx38655, A0=>nx13388, A1=>nx18502);
   ix27902 : oai21 port map ( Y=>nx27901, A0=>nx38661, A1=>nx42723, B0=>
      nx38663);
   booth_booth_integrtaion_6_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_17, QB=>nx38661, D=>nx27901, CLK=>clk, 
      R=>rst);
   ix38664 : nand03 port map ( Y=>nx38663, A0=>nx42731, A1=>nx13896, A2=>
      nx42727);
   ix13897 : xnor2 port map ( Y=>nx13896, A0=>nx38666, A1=>nx18503);
   ix38667 : aoi22 port map ( Y=>nx38666, A0=>
      booth_booth_integration_output_6_17, A1=>nx13412, B0=>nx13388, B1=>
      nx18502);
   ix13403 : nor02_2x port map ( Y=>nx13402, A0=>data_in(96), A1=>
      data_in(97));
   ix27892 : oai21 port map ( Y=>nx27891, A0=>nx38681, A1=>nx42723, B0=>
      nx38683);
   booth_booth_integrtaion_6_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_18, QB=>nx38681, D=>nx27891, CLK=>clk, 
      R=>rst);
   ix38684 : nand03 port map ( Y=>nx38683, A0=>nx42731, A1=>nx13884, A2=>
      nx42727);
   ix13885 : xnor2 port map ( Y=>nx13884, A0=>nx13440, A1=>nx38696);
   ix13441 : oai22 port map ( Y=>nx13440, A0=>nx38666, A1=>nx38687, B0=>
      nx38681, B1=>nx42735);
   ix38690 : aoi32 port map ( Y=>nx38689, A0=>nx13422, A1=>nx42099, A2=>
      nx38692, B0=>data_in(98), B1=>nx42095);
   ix13423 : oai21 port map ( Y=>nx13422, A0=>data_in(96), A1=>data_in(97), 
      B0=>data_in(98));
   ix27882 : oai21 port map ( Y=>nx27881, A0=>nx38700, A1=>nx42723, B0=>
      nx38702);
   booth_booth_integrtaion_6_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_19, QB=>nx38700, D=>nx27881, CLK=>clk, 
      R=>rst);
   ix38703 : nand03 port map ( Y=>nx38702, A0=>nx42731, A1=>nx13872, A2=>
      nx42727);
   ix13873 : xnor2 port map ( Y=>nx13872, A0=>nx38705, A1=>nx18505);
   ix38706 : aoi22 port map ( Y=>nx38705, A0=>
      booth_booth_integration_output_6_19, A1=>nx13460, B0=>nx13440, B1=>
      nx18504);
   ix13461 : oai32 port map ( Y=>nx13460, A0=>nx38708, A1=>nx38671, A2=>
      nx13450, B0=>nx38711, B1=>nx38676);
   ix13427 : nor03_2x port map ( Y=>nx13426, A0=>data_in(98), A1=>
      data_in(96), A2=>data_in(97));
   ix38712 : inv01 port map ( Y=>nx38711, A=>data_in(99));
   ix13451 : nor04 port map ( Y=>nx13450, A0=>data_in(99), A1=>data_in(98), 
      A2=>data_in(96), A3=>data_in(97));
   ix38720 : xnor2 port map ( Y=>nx38719, A0=>nx13488, A1=>nx18507);
   ix13489 : oai22 port map ( Y=>nx13488, A0=>nx38705, A1=>nx38722, B0=>
      nx38733, B1=>nx42737);
   ix38725 : aoi32 port map ( Y=>nx38724, A0=>nx13470, A1=>nx42099, A2=>
      nx38729, B0=>data_in(100), B1=>nx42095);
   ix13471 : nand02 port map ( Y=>nx13470, A0=>nx38727, A1=>data_in(100));
   ix38730 : nand02 port map ( Y=>nx38729, A0=>nx38731, A1=>nx13450);
   ix38732 : inv01 port map ( Y=>nx38731, A=>data_in(100));
   booth_booth_integrtaion_6_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_20, QB=>nx38733, D=>nx27871, CLK=>clk, 
      R=>rst);
   ix27862 : oai21 port map ( Y=>nx27861, A0=>nx38738, A1=>nx42723, B0=>
      nx38740);
   booth_booth_integrtaion_6_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_21, QB=>nx38738, D=>nx27861, CLK=>clk, 
      R=>rst);
   ix38741 : nand03 port map ( Y=>nx38740, A0=>nx42731, A1=>nx13848, A2=>
      nx42727);
   ix13849 : xnor2 port map ( Y=>nx13848, A0=>nx38743, A1=>nx18508);
   ix38744 : aoi22 port map ( Y=>nx38743, A0=>
      booth_booth_integration_output_6_21, A1=>nx13508, B0=>nx13488, B1=>
      nx18507);
   ix13499 : nor02_2x port map ( Y=>nx13498, A0=>data_in(101), A1=>nx38729);
   ix38756 : xnor2 port map ( Y=>nx38755, A0=>nx13536, A1=>nx18509);
   ix13537 : oai22 port map ( Y=>nx13536, A0=>nx38743, A1=>nx38758, B0=>
      nx38769, B1=>nx42739);
   ix38761 : aoi32 port map ( Y=>nx38760, A0=>nx13518, A1=>nx42099, A2=>
      nx38765, B0=>data_in(102), B1=>nx42095);
   ix13519 : nand02 port map ( Y=>nx13518, A0=>nx38763, A1=>data_in(102));
   ix38766 : nand02 port map ( Y=>nx38765, A0=>nx38767, A1=>nx13498);
   ix38768 : inv01 port map ( Y=>nx38767, A=>data_in(102));
   booth_booth_integrtaion_6_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_22, QB=>nx38769, D=>nx27851, CLK=>clk, 
      R=>rst);
   ix27842 : oai21 port map ( Y=>nx27841, A0=>nx38774, A1=>nx42725, B0=>
      nx38776);
   booth_booth_integrtaion_6_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_23, QB=>nx38774, D=>nx27841, CLK=>clk, 
      R=>rst);
   ix38777 : nand03 port map ( Y=>nx38776, A0=>nx42731, A1=>nx13824, A2=>
      nx42727);
   ix13825 : xnor2 port map ( Y=>nx13824, A0=>nx38779, A1=>nx18510);
   ix38780 : aoi22 port map ( Y=>nx38779, A0=>
      booth_booth_integration_output_6_23, A1=>nx13556, B0=>nx13536, B1=>
      nx18509);
   ix13547 : nor02_2x port map ( Y=>nx13546, A0=>data_in(103), A1=>nx38765);
   ix38792 : xnor2 port map ( Y=>nx38791, A0=>nx13584, A1=>nx18511);
   ix13585 : oai22 port map ( Y=>nx13584, A0=>nx38779, A1=>nx38794, B0=>
      nx38805, B1=>nx42741);
   ix38797 : aoi32 port map ( Y=>nx38796, A0=>nx13566, A1=>nx42099, A2=>
      nx38801, B0=>data_in(104), B1=>nx42095);
   ix13567 : nand02 port map ( Y=>nx13566, A0=>nx38799, A1=>data_in(104));
   ix38802 : nand02 port map ( Y=>nx38801, A0=>nx38803, A1=>nx13546);
   ix38804 : inv01 port map ( Y=>nx38803, A=>data_in(104));
   booth_booth_integrtaion_6_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_24, QB=>nx38805, D=>nx27831, CLK=>clk, 
      R=>rst);
   ix27822 : oai21 port map ( Y=>nx27821, A0=>nx38810, A1=>nx42725, B0=>
      nx38812);
   booth_booth_integrtaion_6_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_25, QB=>nx38810, D=>nx27821, CLK=>clk, 
      R=>rst);
   ix38813 : nand03 port map ( Y=>nx38812, A0=>nx42731, A1=>nx13800, A2=>
      nx42727);
   ix13801 : xnor2 port map ( Y=>nx13800, A0=>nx38815, A1=>nx18512);
   ix38816 : aoi22 port map ( Y=>nx38815, A0=>
      booth_booth_integration_output_6_25, A1=>nx13604, B0=>nx13584, B1=>
      nx18511);
   ix13595 : nor02_2x port map ( Y=>nx13594, A0=>data_in(105), A1=>nx38801);
   ix38828 : xnor2 port map ( Y=>nx38827, A0=>nx13632, A1=>nx18513);
   ix13633 : oai22 port map ( Y=>nx13632, A0=>nx38815, A1=>nx38830, B0=>
      nx38841, B1=>nx42743);
   ix38833 : aoi32 port map ( Y=>nx38832, A0=>nx13614, A1=>nx42099, A2=>
      nx38837, B0=>data_in(106), B1=>nx42095);
   ix13615 : nand02 port map ( Y=>nx13614, A0=>nx38835, A1=>data_in(106));
   ix38838 : nand02 port map ( Y=>nx38837, A0=>nx38839, A1=>nx13594);
   ix38840 : inv01 port map ( Y=>nx38839, A=>data_in(106));
   booth_booth_integrtaion_6_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_26, QB=>nx38841, D=>nx27811, CLK=>clk, 
      R=>rst);
   ix27802 : oai21 port map ( Y=>nx27801, A0=>nx38846, A1=>nx42725, B0=>
      nx38848);
   booth_booth_integrtaion_6_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_27, QB=>nx38846, D=>nx27801, CLK=>clk, 
      R=>rst);
   ix38849 : nand03 port map ( Y=>nx38848, A0=>nx43313, A1=>nx13776, A2=>
      nx42727);
   ix13777 : xnor2 port map ( Y=>nx13776, A0=>nx38851, A1=>nx18515);
   ix38852 : aoi22 port map ( Y=>nx38851, A0=>
      booth_booth_integration_output_6_27, A1=>nx13652, B0=>nx13632, B1=>
      nx18513);
   ix13643 : nor02_2x port map ( Y=>nx13642, A0=>data_in(107), A1=>nx38837);
   ix38864 : xnor2 port map ( Y=>nx38863, A0=>nx13680, A1=>nx18517);
   ix13681 : oai22 port map ( Y=>nx13680, A0=>nx38851, A1=>nx38866, B0=>
      nx38877, B1=>nx42745);
   ix38869 : aoi32 port map ( Y=>nx38868, A0=>nx13662, A1=>nx42101, A2=>
      nx38873, B0=>data_in(108), B1=>nx42095);
   ix13663 : nand02 port map ( Y=>nx13662, A0=>nx38871, A1=>data_in(108));
   ix38874 : nand02 port map ( Y=>nx38873, A0=>nx38875, A1=>nx13642);
   ix38876 : inv01 port map ( Y=>nx38875, A=>data_in(108));
   booth_booth_integrtaion_6_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12213, QB=>nx38877, D=>nx27791, CLK=>clk, R=>rst);
   ix27782 : oai21 port map ( Y=>nx27781, A0=>nx38882, A1=>nx42725, B0=>
      nx38884);
   booth_booth_integrtaion_6_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12212, QB=>nx38882, D=>nx27781, CLK=>clk, R=>rst);
   ix38885 : nand03 port map ( Y=>nx38884, A0=>nx43313, A1=>nx13752, A2=>
      nx42725);
   ix13753 : xnor2 port map ( Y=>nx13752, A0=>nx38887, A1=>nx18519);
   ix38888 : aoi22 port map ( Y=>nx38887, A0=>booth_output_29_dup_12212, A1
      =>nx13700, B0=>nx13680, B1=>nx18517);
   ix13691 : nor02_2x port map ( Y=>nx13690, A0=>data_in(109), A1=>nx38873);
   ix27772 : oai21 port map ( Y=>nx27771, A0=>nx38898, A1=>nx42725, B0=>
      nx38900);
   booth_booth_integrtaion_6_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx38898, D=>nx27771, CLK=>clk, R=>rst);
   ix38901 : nand03 port map ( Y=>nx38900, A0=>nx43313, A1=>nx13740, A2=>
      nx42725);
   ix13741 : xnor2 port map ( Y=>nx13740, A0=>nx13728, A1=>nx38915);
   ix13729 : oai22 port map ( Y=>nx13728, A0=>nx38887, A1=>nx38904, B0=>
      nx38898, B1=>nx42747);
   ix38907 : aoi32 port map ( Y=>nx38906, A0=>nx13710, A1=>nx42101, A2=>
      nx38911, B0=>data_in(110), B1=>nx42097);
   ix13711 : nand02 port map ( Y=>nx13710, A0=>nx38909, A1=>data_in(110));
   ix38912 : nand02 port map ( Y=>nx38911, A0=>nx38913, A1=>nx13690);
   ix38914 : inv01 port map ( Y=>nx38913, A=>data_in(110));
   ix13737 : oai22 port map ( Y=>nx13736, A0=>nx38671, A1=>nx38918, B0=>
      nx38920, B1=>nx38676);
   ix38919 : xnor2 port map ( Y=>nx38918, A0=>data_in(111), A1=>nx38911);
   ix38921 : inv01 port map ( Y=>nx38920, A=>data_in(111));
   ix38923 : aoi32 port map ( Y=>nx38922, A0=>nx13686, A1=>nx42101, A2=>
      nx38909, B0=>data_in(109), B1=>nx42097);
   ix13687 : nand02 port map ( Y=>nx13686, A0=>nx38873, A1=>data_in(109));
   ix38926 : aoi32 port map ( Y=>nx38925, A0=>nx13638, A1=>nx42101, A2=>
      nx38871, B0=>data_in(107), B1=>nx42097);
   ix13639 : nand02 port map ( Y=>nx13638, A0=>nx38837, A1=>data_in(107));
   ix38929 : aoi32 port map ( Y=>nx38928, A0=>nx13590, A1=>nx42101, A2=>
      nx38835, B0=>data_in(105), B1=>nx42097);
   ix13591 : nand02 port map ( Y=>nx13590, A0=>nx38801, A1=>data_in(105));
   ix38932 : aoi32 port map ( Y=>nx38931, A0=>nx13542, A1=>nx42101, A2=>
      nx38799, B0=>data_in(103), B1=>nx42097);
   ix13543 : nand02 port map ( Y=>nx13542, A0=>nx38765, A1=>data_in(103));
   ix38935 : aoi32 port map ( Y=>nx38934, A0=>nx13494, A1=>nx42103, A2=>
      nx38763, B0=>data_in(101), B1=>nx42097);
   ix13495 : nand02 port map ( Y=>nx13494, A0=>nx38729, A1=>data_in(101));
   ix38938 : aoi32 port map ( Y=>nx38937, A0=>nx13396, A1=>nx42103, A2=>
      nx38940, B0=>data_in(97), B1=>nx42097);
   ix13397 : nand02 port map ( Y=>nx13396, A0=>data_in(97), A1=>data_in(96)
   );
   booth_booth_integrtaion_6_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_16, QB=>nx38651, D=>nx27911, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_15, QB=>nx38944, D=>nx27921, CLK=>clk, 
      R=>rst);
   ix13977 : aoi21 port map ( Y=>nx13976, A0=>label_7_output_0, A1=>
      booth_booth_integration_output_6_12, B0=>nx43055);
   labelsregfile_label7_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_7_output_1, QB=>nx38961, D=>nx27991, CLK=>clk, R=>rst);
   lat_label_7_input_1 : latch port map ( Q=>label_7_input_1, D=>nx14014, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_1 : dffr port map ( Q=>
      label_7_input_state_machine_1, QB=>OPEN, D=>nx27981, CLK=>clk, R=>rst
   );
   ix14011 : xor2 port map ( Y=>nx14010, A0=>nx38502, A1=>nx38951);
   ix38963 : xnor2 port map ( Y=>nx38962, A0=>
      booth_booth_integration_output_6_14, A1=>label_7_output_2);
   labelsregfile_label7_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_7_output_3, QB=>nx38976, D=>nx28031, CLK=>clk, R=>rst);
   lat_label_7_input_3 : latch port map ( Q=>label_7_input_3, D=>nx14078, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_3 : dffr port map ( Q=>
      label_7_input_state_machine_3, QB=>OPEN, D=>nx28021, CLK=>clk, R=>rst
   );
   ix14075 : xor2 port map ( Y=>nx14074, A0=>nx38491, A1=>nx38966);
   labelsregfile_label7_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_7_output_5, QB=>nx38991, D=>nx28071, CLK=>clk, R=>rst);
   lat_label_7_input_5 : latch port map ( Q=>label_7_input_5, D=>nx14142, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_5 : dffr port map ( Q=>
      label_7_input_state_machine_5, QB=>OPEN, D=>nx28061, CLK=>clk, R=>rst
   );
   ix14139 : xor2 port map ( Y=>nx14138, A0=>nx38480, A1=>nx38981);
   labelsregfile_label7_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_7_output_7, QB=>nx39006, D=>nx28111, CLK=>clk, R=>rst);
   lat_label_7_input_7 : latch port map ( Q=>label_7_input_7, D=>nx14206, 
      CLK=>nx41697);
   reg_label_7_input_state_machine_7 : dffr port map ( Q=>
      label_7_input_state_machine_7, QB=>OPEN, D=>nx28101, CLK=>clk, R=>rst
   );
   ix14203 : xor2 port map ( Y=>nx14202, A0=>nx38469, A1=>nx38996);
   labelsregfile_label7_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_7_output_9, QB=>nx39021, D=>nx28151, CLK=>clk, R=>rst);
   lat_label_7_input_9 : latch port map ( Q=>label_7_input_9, D=>nx14270, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_9 : dffr port map ( Q=>
      label_7_input_state_machine_9, QB=>OPEN, D=>nx28141, CLK=>clk, R=>rst
   );
   ix14267 : xor2 port map ( Y=>nx14266, A0=>nx38458, A1=>nx39011);
   labelsregfile_label7_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_7_output_11, QB=>nx39036, D=>nx28191, CLK=>clk, R=>rst);
   lat_label_7_input_11 : latch port map ( Q=>label_7_input_11, D=>nx14334, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_11 : dffr port map ( Q=>
      label_7_input_state_machine_11, QB=>OPEN, D=>nx28181, CLK=>clk, R=>rst
   );
   ix14331 : xor2 port map ( Y=>nx14330, A0=>nx38447, A1=>nx39026);
   labelsregfile_label7_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_7_output_13, QB=>nx39051, D=>nx28231, CLK=>clk, R=>rst);
   lat_label_7_input_13 : latch port map ( Q=>label_7_input_13, D=>nx14398, 
      CLK=>nx41699);
   reg_label_7_input_state_machine_13 : dffr port map ( Q=>
      label_7_input_state_machine_13, QB=>OPEN, D=>nx28221, CLK=>clk, R=>rst
   );
   ix14395 : xor2 port map ( Y=>nx14394, A0=>nx38436, A1=>nx39041);
   ix29092 : oai21 port map ( Y=>nx29091, A0=>nx39057, A1=>nx41625, B0=>
      nx39059);
   max_calc_reg_comparator_fourth_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx39057, D=>nx29091, CLK=>clk);
   ix39060 : nand03 port map ( Y=>nx39059, A0=>label_8_output_14, A1=>
      nx42639, A2=>nx41625);
   labelsregfile_label8_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_8_output_14, QB=>OPEN, D=>nx29081, CLK=>clk, R=>rst);
   lat_label_8_input_14 : latch port map ( Q=>label_8_input_14, D=>nx15740, 
      CLK=>nx41705);
   reg_label_8_input_state_machine_14 : dffr port map ( Q=>
      label_8_input_state_machine_14, QB=>OPEN, D=>nx28261, CLK=>clk, R=>rst
   );
   ix15737 : xnor2 port map ( Y=>nx15736, A0=>nx15732, A1=>nx39686);
   ix15733 : oai22 port map ( Y=>nx15732, A0=>nx39070, A1=>nx39675, B0=>
      nx39685, B1=>nx39444);
   ix39071 : aoi22 port map ( Y=>nx39070, A0=>label_8_output_12, A1=>
      booth_booth_integration_output_7_24, B0=>nx15668, B1=>nx18580);
   labelsregfile_label8_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_8_output_12, QB=>OPEN, D=>nx29051, CLK=>clk, R=>rst);
   lat_label_8_input_12 : latch port map ( Q=>label_8_input_12, D=>nx15682, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_12 : dffr port map ( Q=>
      label_8_input_state_machine_12, QB=>OPEN, D=>nx29041, CLK=>clk, R=>rst
   );
   ix15679 : xnor2 port map ( Y=>nx15678, A0=>nx15668, A1=>nx39671);
   ix15669 : oai22 port map ( Y=>nx15668, A0=>nx39081, A1=>nx39660, B0=>
      nx39670, B1=>nx39408);
   ix39082 : aoi22 port map ( Y=>nx39081, A0=>label_8_output_10, A1=>
      booth_booth_integration_output_7_22, B0=>nx15604, B1=>nx18578);
   labelsregfile_label8_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_8_output_10, QB=>OPEN, D=>nx29011, CLK=>clk, R=>rst);
   lat_label_8_input_10 : latch port map ( Q=>label_8_input_10, D=>nx15618, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_10 : dffr port map ( Q=>
      label_8_input_state_machine_10, QB=>OPEN, D=>nx29001, CLK=>clk, R=>rst
   );
   ix15615 : xnor2 port map ( Y=>nx15614, A0=>nx15604, A1=>nx39656);
   ix15605 : oai22 port map ( Y=>nx15604, A0=>nx39092, A1=>nx39645, B0=>
      nx39655, B1=>nx39372);
   ix39093 : aoi22 port map ( Y=>nx39092, A0=>label_8_output_8, A1=>
      booth_booth_integration_output_7_20, B0=>nx15540, B1=>nx18576);
   labelsregfile_label8_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_8_output_8, QB=>OPEN, D=>nx28971, CLK=>clk, R=>rst);
   lat_label_8_input_8 : latch port map ( Q=>label_8_input_8, D=>nx15554, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_8 : dffr port map ( Q=>
      label_8_input_state_machine_8, QB=>OPEN, D=>nx28961, CLK=>clk, R=>rst
   );
   ix15551 : xnor2 port map ( Y=>nx15550, A0=>nx15540, A1=>nx39641);
   ix15541 : oai22 port map ( Y=>nx15540, A0=>nx39103, A1=>nx39630, B0=>
      nx39640, B1=>nx39334);
   ix39104 : aoi22 port map ( Y=>nx39103, A0=>label_8_output_6, A1=>
      booth_booth_integration_output_7_18, B0=>nx15476, B1=>nx18573);
   labelsregfile_label8_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_8_output_6, QB=>OPEN, D=>nx28931, CLK=>clk, R=>rst);
   lat_label_8_input_6 : latch port map ( Q=>label_8_input_6, D=>nx15490, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_6 : dffr port map ( Q=>
      label_8_input_state_machine_6, QB=>OPEN, D=>nx28921, CLK=>clk, R=>rst
   );
   ix15487 : xnor2 port map ( Y=>nx15486, A0=>nx15476, A1=>nx39626);
   ix15477 : oai22 port map ( Y=>nx15476, A0=>nx39114, A1=>nx39615, B0=>
      nx39625, B1=>nx39295);
   ix39115 : aoi22 port map ( Y=>nx39114, A0=>label_8_output_4, A1=>
      booth_booth_integration_output_7_16, B0=>nx15412, B1=>nx18569);
   labelsregfile_label8_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_8_output_4, QB=>OPEN, D=>nx28891, CLK=>clk, R=>rst);
   lat_label_8_input_4 : latch port map ( Q=>label_8_input_4, D=>nx15426, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_4 : dffr port map ( Q=>
      label_8_input_state_machine_4, QB=>OPEN, D=>nx28881, CLK=>clk, R=>rst
   );
   ix15423 : xnor2 port map ( Y=>nx15422, A0=>nx15412, A1=>nx39611);
   ix15413 : oai22 port map ( Y=>nx15412, A0=>nx39125, A1=>nx39600, B0=>
      nx39610, B1=>nx39578);
   ix39126 : aoi22 port map ( Y=>nx39125, A0=>label_8_output_2, A1=>
      booth_booth_integration_output_7_14, B0=>nx15348, B1=>nx18566);
   labelsregfile_label8_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_8_output_2, QB=>OPEN, D=>nx28851, CLK=>clk, R=>rst);
   lat_label_8_input_2 : latch port map ( Q=>label_8_input_2, D=>nx15362, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_2 : dffr port map ( Q=>
      label_8_input_state_machine_2, QB=>OPEN, D=>nx28841, CLK=>clk, R=>rst
   );
   ix15359 : xnor2 port map ( Y=>nx15358, A0=>nx15348, A1=>nx39596);
   ix15349 : oai22 port map ( Y=>nx15348, A0=>nx39136, A1=>nx39585, B0=>
      nx39595, B1=>nx39581);
   ix39137 : nand02 port map ( Y=>nx39136, A0=>label_8_output_0, A1=>
      booth_booth_integration_output_7_12);
   labelsregfile_label8_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_8_output_0, QB=>OPEN, D=>nx28811, CLK=>clk, R=>rst);
   lat_label_8_input_0 : latch port map ( Q=>label_8_input_0, D=>nx15304, 
      CLK=>nx41701);
   ix15305 : oai21 port map ( Y=>nx15304, A0=>nx39142, A1=>nx41461, B0=>
      nx39146);
   reg_label_8_input_state_machine_0 : dffr port map ( Q=>
      label_8_input_state_machine_0, QB=>nx39142, D=>nx28801, CLK=>clk, R=>
      rst);
   ix39147 : oai21 port map ( Y=>nx39146, A0=>
      booth_booth_integration_output_7_12, A1=>label_8_output_0, B0=>nx15292
   );
   booth_booth_integrtaion_7_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_12, QB=>OPEN, D=>nx28791, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_13, QB=>nx39581, D=>nx28781, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_14, QB=>OPEN, D=>nx28771, CLK=>clk, R
      =>rst);
   ix39160 : aoi22 port map ( Y=>nx39159, A0=>nx41797, A1=>nx42119, B0=>
      nx15234, B1=>nx15240);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_reg_output_0, QB=>OPEN, 
      D=>nx28291, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_0, QB=>OPEN, D=>nx28277, CLK
      =>clk, S=>nx41505);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_reg_output_9, QB=>OPEN, 
      D=>nx28471, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_9, QB=>OPEN, D=>nx28461, CLK
      =>clk, R=>nx41505);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>output_8_dup_12884, QB=>OPEN, D=>nx28451, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_8, QB=>OPEN, D=>nx28441, CLK
      =>clk, R=>nx41505);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>output_7_dup_12885, QB=>OPEN, D=>nx28431, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_7, QB=>OPEN, D=>nx28421, CLK
      =>clk, R=>nx41505);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>output_6_dup_12886, QB=>OPEN, D=>nx28411, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_6, QB=>OPEN, D=>nx28401, CLK
      =>clk, R=>nx41505);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>output_5_dup_12887, QB=>OPEN, D=>nx28391, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_5, QB=>OPEN, D=>nx28381, CLK
      =>clk, R=>nx41503);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>output_4_dup_12888, QB=>OPEN, D=>nx28371, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_4, QB=>OPEN, D=>nx28361, CLK
      =>clk, R=>nx41503);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>output_3_dup_12889, QB=>OPEN, D=>nx28351, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_3, QB=>OPEN, D=>nx28341, CLK
      =>clk, R=>nx41503);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>output_2_dup_12890, QB=>OPEN, D=>nx28331, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_2, QB=>OPEN, D=>nx28321, CLK
      =>clk, R=>nx41503);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>output_1_dup_12891, QB=>OPEN, D=>nx28311, CLK=>clk, R=>
      rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_1, QB=>OPEN, D=>nx28301, CLK
      =>clk, R=>nx41503);
   ix28272 : nand02 port map ( Y=>nx28271, A0=>nx42961, A1=>nx42105);
   booth_booth_integrtaion_7_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx39206, D=>nx28271, CLK=>clk, S=>nx41503);
   ix15235 : nand02 port map ( Y=>nx15234, A0=>nx39227, A1=>nx39285);
   ix39228 : oai21 port map ( Y=>nx39227, A0=>nx42131, A1=>nx42127, B0=>
      data_in(112));
   ix28602 : oai21 port map ( Y=>nx28601, A0=>nx39232, A1=>nx42749, B0=>
      nx39234);
   booth_booth_integrtaion_7_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx39232, D=>nx28601, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_output_0_dup_12244, QB=>nx39283, D=>nx28591, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_output_1_dup_12243, QB=>OPEN, D=>nx28581, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_output_2_dup_12242, QB=>OPEN, D=>nx28571, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_output_3_dup_12241, QB=>OPEN, D=>nx28561, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_output_4_dup_12240, QB=>OPEN, D=>nx28551, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_output_5_dup_12239, QB=>OPEN, D=>nx28541, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_output_6_dup_12238, QB=>OPEN, D=>nx28531, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_output_7_dup_12237, QB=>OPEN, D=>nx28521, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_output_8_dup_12236, QB=>OPEN, D=>nx28511, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_output_9_dup_12235, QB=>OPEN, D=>nx28501, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_output_10_dup_12234, QB=>OPEN, D=>nx28491, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_output_11_dup_12233, QB=>OPEN, D=>nx28481, CLK=>clk, R=>rst);
   ix39290 : xnor2 port map ( Y=>nx39289, A0=>nx14704, A1=>nx18544);
   ix28742 : oai21 port map ( Y=>nx28741, A0=>nx39295, A1=>nx42749, B0=>
      nx39297);
   booth_booth_integrtaion_7_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_17, QB=>nx39295, D=>nx28741, CLK=>clk, 
      R=>rst);
   ix39298 : nand03 port map ( Y=>nx39297, A0=>nx42757, A1=>nx15212, A2=>
      nx42753);
   ix15213 : xnor2 port map ( Y=>nx15212, A0=>nx39300, A1=>nx18545);
   ix39301 : aoi22 port map ( Y=>nx39300, A0=>
      booth_booth_integration_output_7_17, A1=>nx14728, B0=>nx14704, B1=>
      nx18544);
   ix14719 : nor02_2x port map ( Y=>nx14718, A0=>data_in(112), A1=>
      data_in(113));
   ix28732 : oai21 port map ( Y=>nx28731, A0=>nx39315, A1=>nx42749, B0=>
      nx39317);
   booth_booth_integrtaion_7_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_18, QB=>nx39315, D=>nx28731, CLK=>clk, 
      R=>rst);
   ix39318 : nand03 port map ( Y=>nx39317, A0=>nx42757, A1=>nx15200, A2=>
      nx42753);
   ix15201 : xnor2 port map ( Y=>nx15200, A0=>nx14756, A1=>nx39330);
   ix14757 : oai22 port map ( Y=>nx14756, A0=>nx39300, A1=>nx39321, B0=>
      nx39315, B1=>nx42761);
   ix39324 : aoi32 port map ( Y=>nx39323, A0=>nx14738, A1=>nx42131, A2=>
      nx39326, B0=>data_in(114), B1=>nx42127);
   ix14739 : oai21 port map ( Y=>nx14738, A0=>data_in(112), A1=>data_in(113), 
      B0=>data_in(114));
   ix28722 : oai21 port map ( Y=>nx28721, A0=>nx39334, A1=>nx42749, B0=>
      nx39336);
   booth_booth_integrtaion_7_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_19, QB=>nx39334, D=>nx28721, CLK=>clk, 
      R=>rst);
   ix39337 : nand03 port map ( Y=>nx39336, A0=>nx42757, A1=>nx15188, A2=>
      nx42753);
   ix15189 : xnor2 port map ( Y=>nx15188, A0=>nx39339, A1=>nx18547);
   ix39340 : aoi22 port map ( Y=>nx39339, A0=>
      booth_booth_integration_output_7_19, A1=>nx14776, B0=>nx14756, B1=>
      nx18546);
   ix14777 : oai32 port map ( Y=>nx14776, A0=>nx39342, A1=>nx39305, A2=>
      nx14766, B0=>nx39345, B1=>nx39310);
   ix14743 : nor03_2x port map ( Y=>nx14742, A0=>data_in(114), A1=>
      data_in(112), A2=>data_in(113));
   ix39346 : inv01 port map ( Y=>nx39345, A=>data_in(115));
   ix14767 : nor04 port map ( Y=>nx14766, A0=>data_in(115), A1=>data_in(114), 
      A2=>data_in(112), A3=>data_in(113));
   ix39354 : xnor2 port map ( Y=>nx39353, A0=>nx14804, A1=>nx18548);
   ix14805 : oai22 port map ( Y=>nx14804, A0=>nx39339, A1=>nx39356, B0=>
      nx39367, B1=>nx42763);
   ix39359 : aoi32 port map ( Y=>nx39358, A0=>nx14786, A1=>nx42131, A2=>
      nx39363, B0=>data_in(116), B1=>nx42127);
   ix14787 : nand02 port map ( Y=>nx14786, A0=>nx39361, A1=>data_in(116));
   ix39364 : nand02 port map ( Y=>nx39363, A0=>nx39365, A1=>nx14766);
   ix39366 : inv01 port map ( Y=>nx39365, A=>data_in(116));
   booth_booth_integrtaion_7_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_20, QB=>nx39367, D=>nx28711, CLK=>clk, 
      R=>rst);
   ix28702 : oai21 port map ( Y=>nx28701, A0=>nx39372, A1=>nx42749, B0=>
      nx39374);
   booth_booth_integrtaion_7_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_21, QB=>nx39372, D=>nx28701, CLK=>clk, 
      R=>rst);
   ix39375 : nand03 port map ( Y=>nx39374, A0=>nx42757, A1=>nx15164, A2=>
      nx42753);
   ix15165 : xnor2 port map ( Y=>nx15164, A0=>nx39377, A1=>nx18549);
   ix39378 : aoi22 port map ( Y=>nx39377, A0=>
      booth_booth_integration_output_7_21, A1=>nx14824, B0=>nx14804, B1=>
      nx18548);
   ix14815 : nor02_2x port map ( Y=>nx14814, A0=>data_in(117), A1=>nx39363);
   ix39390 : xnor2 port map ( Y=>nx39389, A0=>nx14852, A1=>nx18551);
   ix14853 : oai22 port map ( Y=>nx14852, A0=>nx39377, A1=>nx39392, B0=>
      nx39403, B1=>nx42765);
   ix39395 : aoi32 port map ( Y=>nx39394, A0=>nx14834, A1=>nx42131, A2=>
      nx39399, B0=>data_in(118), B1=>nx42127);
   ix14835 : nand02 port map ( Y=>nx14834, A0=>nx39397, A1=>data_in(118));
   ix39400 : nand02 port map ( Y=>nx39399, A0=>nx39401, A1=>nx14814);
   ix39402 : inv01 port map ( Y=>nx39401, A=>data_in(118));
   booth_booth_integrtaion_7_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_22, QB=>nx39403, D=>nx28691, CLK=>clk, 
      R=>rst);
   ix28682 : oai21 port map ( Y=>nx28681, A0=>nx39408, A1=>nx42751, B0=>
      nx39410);
   booth_booth_integrtaion_7_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_23, QB=>nx39408, D=>nx28681, CLK=>clk, 
      R=>rst);
   ix39411 : nand03 port map ( Y=>nx39410, A0=>nx42757, A1=>nx15140, A2=>
      nx42753);
   ix15141 : xnor2 port map ( Y=>nx15140, A0=>nx39413, A1=>nx18553);
   ix39414 : aoi22 port map ( Y=>nx39413, A0=>
      booth_booth_integration_output_7_23, A1=>nx14872, B0=>nx14852, B1=>
      nx18551);
   ix14863 : nor02_2x port map ( Y=>nx14862, A0=>data_in(119), A1=>nx39399);
   ix39426 : xnor2 port map ( Y=>nx39425, A0=>nx14900, A1=>nx18555);
   ix14901 : oai22 port map ( Y=>nx14900, A0=>nx39413, A1=>nx39428, B0=>
      nx39439, B1=>nx42767);
   ix39431 : aoi32 port map ( Y=>nx39430, A0=>nx14882, A1=>nx42131, A2=>
      nx39435, B0=>data_in(120), B1=>nx42127);
   ix14883 : nand02 port map ( Y=>nx14882, A0=>nx39433, A1=>data_in(120));
   ix39436 : nand02 port map ( Y=>nx39435, A0=>nx39437, A1=>nx14862);
   ix39438 : inv01 port map ( Y=>nx39437, A=>data_in(120));
   booth_booth_integrtaion_7_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_24, QB=>nx39439, D=>nx28671, CLK=>clk, 
      R=>rst);
   ix28662 : oai21 port map ( Y=>nx28661, A0=>nx39444, A1=>nx42751, B0=>
      nx39446);
   booth_booth_integrtaion_7_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_25, QB=>nx39444, D=>nx28661, CLK=>clk, 
      R=>rst);
   ix39447 : nand03 port map ( Y=>nx39446, A0=>nx42757, A1=>nx15116, A2=>
      nx42753);
   ix15117 : xnor2 port map ( Y=>nx15116, A0=>nx39449, A1=>nx18557);
   ix39450 : aoi22 port map ( Y=>nx39449, A0=>
      booth_booth_integration_output_7_25, A1=>nx14920, B0=>nx14900, B1=>
      nx18555);
   ix14911 : nor02_2x port map ( Y=>nx14910, A0=>data_in(121), A1=>nx39435);
   ix39462 : xnor2 port map ( Y=>nx39461, A0=>nx14948, A1=>nx18559);
   ix14949 : oai22 port map ( Y=>nx14948, A0=>nx39449, A1=>nx39464, B0=>
      nx39475, B1=>nx42769);
   ix39467 : aoi32 port map ( Y=>nx39466, A0=>nx14930, A1=>nx42131, A2=>
      nx39471, B0=>data_in(122), B1=>nx42127);
   ix14931 : nand02 port map ( Y=>nx14930, A0=>nx39469, A1=>data_in(122));
   ix39472 : nand02 port map ( Y=>nx39471, A0=>nx39473, A1=>nx14910);
   ix39474 : inv01 port map ( Y=>nx39473, A=>data_in(122));
   booth_booth_integrtaion_7_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_26, QB=>nx39475, D=>nx28651, CLK=>clk, 
      R=>rst);
   ix28642 : oai21 port map ( Y=>nx28641, A0=>nx39480, A1=>nx42751, B0=>
      nx39482);
   booth_booth_integrtaion_7_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_27, QB=>nx39480, D=>nx28641, CLK=>clk, 
      R=>rst);
   ix39483 : nand03 port map ( Y=>nx39482, A0=>nx43327, A1=>nx15092, A2=>
      nx42753);
   ix15093 : xnor2 port map ( Y=>nx15092, A0=>nx39485, A1=>nx18561);
   ix39486 : aoi22 port map ( Y=>nx39485, A0=>
      booth_booth_integration_output_7_27, A1=>nx14968, B0=>nx14948, B1=>
      nx18559);
   ix14959 : nor02_2x port map ( Y=>nx14958, A0=>data_in(123), A1=>nx39471);
   ix39498 : xnor2 port map ( Y=>nx39497, A0=>nx14996, A1=>nx18562);
   ix14997 : oai22 port map ( Y=>nx14996, A0=>nx39485, A1=>nx39500, B0=>
      nx39511, B1=>nx42771);
   ix39503 : aoi32 port map ( Y=>nx39502, A0=>nx14978, A1=>nx42133, A2=>
      nx39507, B0=>data_in(124), B1=>nx42127);
   ix14979 : nand02 port map ( Y=>nx14978, A0=>nx39505, A1=>data_in(124));
   ix39508 : nand02 port map ( Y=>nx39507, A0=>nx39509, A1=>nx14958);
   ix39510 : inv01 port map ( Y=>nx39509, A=>data_in(124));
   booth_booth_integrtaion_7_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_output_28_dup_12232, QB=>nx39511, D=>nx28631, CLK=>clk, R=>rst);
   ix28622 : oai21 port map ( Y=>nx28621, A0=>nx39516, A1=>nx42751, B0=>
      nx39518);
   booth_booth_integrtaion_7_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_output_29_dup_12231, QB=>nx39516, D=>nx28621, CLK=>clk, R=>rst);
   ix39519 : nand03 port map ( Y=>nx39518, A0=>nx43327, A1=>nx15068, A2=>
      nx42751);
   ix15069 : xnor2 port map ( Y=>nx15068, A0=>nx39521, A1=>nx18563);
   ix39522 : aoi22 port map ( Y=>nx39521, A0=>booth_output_29_dup_12231, A1
      =>nx15016, B0=>nx14996, B1=>nx18562);
   ix15007 : nor02_2x port map ( Y=>nx15006, A0=>data_in(125), A1=>nx39507);
   ix28612 : oai21 port map ( Y=>nx28611, A0=>nx39532, A1=>nx42751, B0=>
      nx39534);
   booth_booth_integrtaion_7_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx39532, D=>nx28611, CLK=>clk, R=>rst);
   ix39535 : nand03 port map ( Y=>nx39534, A0=>nx43327, A1=>nx15056, A2=>
      nx42751);
   ix15057 : xnor2 port map ( Y=>nx15056, A0=>nx15044, A1=>nx39549);
   ix15045 : oai22 port map ( Y=>nx15044, A0=>nx39521, A1=>nx39538, B0=>
      nx39532, B1=>nx42773);
   ix39541 : aoi32 port map ( Y=>nx39540, A0=>nx15026, A1=>nx42133, A2=>
      nx39545, B0=>data_in(126), B1=>nx42129);
   ix15027 : nand02 port map ( Y=>nx15026, A0=>nx39543, A1=>data_in(126));
   ix39546 : nand02 port map ( Y=>nx39545, A0=>nx39547, A1=>nx15006);
   ix39548 : inv01 port map ( Y=>nx39547, A=>data_in(126));
   ix15053 : oai22 port map ( Y=>nx15052, A0=>nx39305, A1=>nx39552, B0=>
      nx39554, B1=>nx39310);
   ix39553 : xnor2 port map ( Y=>nx39552, A0=>data_in(127), A1=>nx39545);
   ix39555 : inv01 port map ( Y=>nx39554, A=>data_in(127));
   ix39557 : aoi32 port map ( Y=>nx39556, A0=>nx15002, A1=>nx42133, A2=>
      nx39543, B0=>data_in(125), B1=>nx42129);
   ix15003 : nand02 port map ( Y=>nx15002, A0=>nx39507, A1=>data_in(125));
   ix39560 : aoi32 port map ( Y=>nx39559, A0=>nx14954, A1=>nx42133, A2=>
      nx39505, B0=>data_in(123), B1=>nx42129);
   ix14955 : nand02 port map ( Y=>nx14954, A0=>nx39471, A1=>data_in(123));
   ix39563 : aoi32 port map ( Y=>nx39562, A0=>nx14906, A1=>nx42133, A2=>
      nx39469, B0=>data_in(121), B1=>nx42129);
   ix14907 : nand02 port map ( Y=>nx14906, A0=>nx39435, A1=>data_in(121));
   ix39566 : aoi32 port map ( Y=>nx39565, A0=>nx14858, A1=>nx42133, A2=>
      nx39433, B0=>data_in(119), B1=>nx42129);
   ix14859 : nand02 port map ( Y=>nx14858, A0=>nx39399, A1=>data_in(119));
   ix39569 : aoi32 port map ( Y=>nx39568, A0=>nx14810, A1=>nx42135, A2=>
      nx39397, B0=>data_in(117), B1=>nx42129);
   ix14811 : nand02 port map ( Y=>nx14810, A0=>nx39363, A1=>data_in(117));
   ix39572 : aoi32 port map ( Y=>nx39571, A0=>nx14712, A1=>nx42135, A2=>
      nx39574, B0=>data_in(113), B1=>nx42129);
   ix14713 : nand02 port map ( Y=>nx14712, A0=>data_in(113), A1=>
      data_in(112));
   booth_booth_integrtaion_7_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_16, QB=>nx39285, D=>nx28751, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_15, QB=>nx39578, D=>nx28761, CLK=>clk, 
      R=>rst);
   ix15293 : aoi21 port map ( Y=>nx15292, A0=>label_8_output_0, A1=>
      booth_booth_integration_output_7_12, B0=>nx43055);
   labelsregfile_label8_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_8_output_1, QB=>nx39595, D=>nx28831, CLK=>clk, R=>rst);
   lat_label_8_input_1 : latch port map ( Q=>label_8_input_1, D=>nx15330, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_1 : dffr port map ( Q=>
      label_8_input_state_machine_1, QB=>OPEN, D=>nx28821, CLK=>clk, R=>rst
   );
   ix15327 : xor2 port map ( Y=>nx15326, A0=>nx39136, A1=>nx39585);
   ix39597 : xnor2 port map ( Y=>nx39596, A0=>
      booth_booth_integration_output_7_14, A1=>label_8_output_2);
   labelsregfile_label8_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_8_output_3, QB=>nx39610, D=>nx28871, CLK=>clk, R=>rst);
   lat_label_8_input_3 : latch port map ( Q=>label_8_input_3, D=>nx15394, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_3 : dffr port map ( Q=>
      label_8_input_state_machine_3, QB=>OPEN, D=>nx28861, CLK=>clk, R=>rst
   );
   ix15391 : xor2 port map ( Y=>nx15390, A0=>nx39125, A1=>nx39600);
   labelsregfile_label8_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_8_output_5, QB=>nx39625, D=>nx28911, CLK=>clk, R=>rst);
   lat_label_8_input_5 : latch port map ( Q=>label_8_input_5, D=>nx15458, 
      CLK=>nx41701);
   reg_label_8_input_state_machine_5 : dffr port map ( Q=>
      label_8_input_state_machine_5, QB=>OPEN, D=>nx28901, CLK=>clk, R=>rst
   );
   ix15455 : xor2 port map ( Y=>nx15454, A0=>nx39114, A1=>nx39615);
   labelsregfile_label8_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_8_output_7, QB=>nx39640, D=>nx28951, CLK=>clk, R=>rst);
   lat_label_8_input_7 : latch port map ( Q=>label_8_input_7, D=>nx15522, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_7 : dffr port map ( Q=>
      label_8_input_state_machine_7, QB=>OPEN, D=>nx28941, CLK=>clk, R=>rst
   );
   ix15519 : xor2 port map ( Y=>nx15518, A0=>nx39103, A1=>nx39630);
   labelsregfile_label8_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_8_output_9, QB=>nx39655, D=>nx28991, CLK=>clk, R=>rst);
   lat_label_8_input_9 : latch port map ( Q=>label_8_input_9, D=>nx15586, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_9 : dffr port map ( Q=>
      label_8_input_state_machine_9, QB=>OPEN, D=>nx28981, CLK=>clk, R=>rst
   );
   ix15583 : xor2 port map ( Y=>nx15582, A0=>nx39092, A1=>nx39645);
   labelsregfile_label8_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_8_output_11, QB=>nx39670, D=>nx29031, CLK=>clk, R=>rst);
   lat_label_8_input_11 : latch port map ( Q=>label_8_input_11, D=>nx15650, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_11 : dffr port map ( Q=>
      label_8_input_state_machine_11, QB=>OPEN, D=>nx29021, CLK=>clk, R=>rst
   );
   ix15647 : xor2 port map ( Y=>nx15646, A0=>nx39081, A1=>nx39660);
   labelsregfile_label8_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_8_output_13, QB=>nx39685, D=>nx29071, CLK=>clk, R=>rst);
   lat_label_8_input_13 : latch port map ( Q=>label_8_input_13, D=>nx15714, 
      CLK=>nx41703);
   reg_label_8_input_state_machine_13 : dffr port map ( Q=>
      label_8_input_state_machine_13, QB=>OPEN, D=>nx29061, CLK=>clk, R=>rst
   );
   ix15711 : xor2 port map ( Y=>nx15710, A0=>nx39070, A1=>nx39675);
   ix16277 : xnor2 port map ( Y=>nx16276, A0=>nx39690, A1=>nx16274);
   ix39691 : aoi22 port map ( Y=>nx39690, A0=>nx39057, A1=>
      max_calc_comparator_fourth_inp1_14, B0=>nx15762, B1=>nx16180);
   ix16181 : oai22 port map ( Y=>nx16180, A0=>nx39694, A1=>nx39707, B0=>
      max_calc_comparator_fourth_inp2_13, B1=>nx39702);
   ix29102 : oai21 port map ( Y=>nx29101, A0=>nx39698, A1=>nx41625, B0=>
      nx39700);
   max_calc_reg_comparator_fourth_inp2_13 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_13, QB=>nx39698, D=>nx29101, CLK=>clk
   );
   max_calc_reg_comparator_fourth_inp1_13 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_13, QB=>nx39702, D=>nx29111, CLK=>clk
   );
   ix29112 : oai21 port map ( Y=>nx29111, A0=>nx39702, A1=>nx41625, B0=>
      nx39705);
   ix39708 : aoi22 port map ( Y=>nx39707, A0=>nx39709, A1=>
      max_calc_comparator_fourth_inp1_12, B0=>nx15806, B1=>nx16164);
   max_calc_reg_comparator_fourth_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx39709, D=>nx29121, CLK=>clk);
   ix29122 : oai21 port map ( Y=>nx29121, A0=>nx39709, A1=>nx41625, B0=>
      nx39712);
   ix39713 : nand03 port map ( Y=>nx39712, A0=>label_8_output_12, A1=>
      nx42641, A2=>nx41627);
   ix29132 : oai21 port map ( Y=>nx29131, A0=>nx39716, A1=>nx41627, B0=>
      nx39718);
   max_calc_reg_comparator_fourth_inp1_12 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_12, QB=>nx39716, D=>nx29131, CLK=>clk
   );
   ix39719 : nand03 port map ( Y=>nx39718, A0=>label_7_output_12, A1=>
      nx42641, A2=>nx41627);
   ix16165 : oai22 port map ( Y=>nx16164, A0=>nx39722, A1=>nx39735, B0=>
      max_calc_comparator_fourth_inp2_11, B1=>nx39730);
   ix29142 : oai21 port map ( Y=>nx29141, A0=>nx39726, A1=>nx41627, B0=>
      nx39728);
   max_calc_reg_comparator_fourth_inp2_11 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_11, QB=>nx39726, D=>nx29141, CLK=>clk
   );
   max_calc_reg_comparator_fourth_inp1_11 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_11, QB=>nx39730, D=>nx29151, CLK=>clk
   );
   ix29152 : oai21 port map ( Y=>nx29151, A0=>nx39730, A1=>nx41627, B0=>
      nx39733);
   ix39736 : aoi22 port map ( Y=>nx39735, A0=>nx39737, A1=>
      max_calc_comparator_fourth_inp1_10, B0=>nx15850, B1=>nx16148);
   max_calc_reg_comparator_fourth_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx39737, D=>nx29161, CLK=>clk);
   ix29162 : oai21 port map ( Y=>nx29161, A0=>nx39737, A1=>nx41629, B0=>
      nx39740);
   ix39741 : nand03 port map ( Y=>nx39740, A0=>label_8_output_10, A1=>
      nx42641, A2=>nx41629);
   ix29172 : oai21 port map ( Y=>nx29171, A0=>nx39744, A1=>nx41629, B0=>
      nx39746);
   max_calc_reg_comparator_fourth_inp1_10 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_10, QB=>nx39744, D=>nx29171, CLK=>clk
   );
   ix39747 : nand03 port map ( Y=>nx39746, A0=>label_7_output_10, A1=>
      nx42641, A2=>nx41629);
   ix16149 : oai22 port map ( Y=>nx16148, A0=>nx39750, A1=>nx39763, B0=>
      max_calc_comparator_fourth_inp2_9, B1=>nx39758);
   ix29182 : oai21 port map ( Y=>nx29181, A0=>nx39754, A1=>nx41629, B0=>
      nx39756);
   max_calc_reg_comparator_fourth_inp2_9 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_9, QB=>nx39754, D=>nx29181, CLK=>clk);
   max_calc_reg_comparator_fourth_inp1_9 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_9, QB=>nx39758, D=>nx29191, CLK=>clk);
   ix29192 : oai21 port map ( Y=>nx29191, A0=>nx39758, A1=>nx41629, B0=>
      nx39761);
   ix39764 : aoi22 port map ( Y=>nx39763, A0=>nx39765, A1=>
      max_calc_comparator_fourth_inp1_8, B0=>nx15894, B1=>nx16132);
   max_calc_reg_comparator_fourth_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx39765, D=>nx29201, CLK=>clk);
   ix29202 : oai21 port map ( Y=>nx29201, A0=>nx39765, A1=>nx41631, B0=>
      nx39768);
   ix39769 : nand03 port map ( Y=>nx39768, A0=>label_8_output_8, A1=>nx42643, 
      A2=>nx41631);
   ix29212 : oai21 port map ( Y=>nx29211, A0=>nx39772, A1=>nx41631, B0=>
      nx39774);
   max_calc_reg_comparator_fourth_inp1_8 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_8, QB=>nx39772, D=>nx29211, CLK=>clk);
   ix39775 : nand03 port map ( Y=>nx39774, A0=>label_7_output_8, A1=>nx42643, 
      A2=>nx41631);
   ix16133 : oai22 port map ( Y=>nx16132, A0=>nx39778, A1=>nx39791, B0=>
      max_calc_comparator_fourth_inp2_7, B1=>nx39786);
   ix29222 : oai21 port map ( Y=>nx29221, A0=>nx39782, A1=>nx41631, B0=>
      nx39784);
   max_calc_reg_comparator_fourth_inp2_7 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_7, QB=>nx39782, D=>nx29221, CLK=>clk);
   max_calc_reg_comparator_fourth_inp1_7 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_7, QB=>nx39786, D=>nx29231, CLK=>clk);
   ix29232 : oai21 port map ( Y=>nx29231, A0=>nx39786, A1=>nx41633, B0=>
      nx39789);
   ix39792 : aoi22 port map ( Y=>nx39791, A0=>nx39793, A1=>
      max_calc_comparator_fourth_inp1_6, B0=>nx15938, B1=>nx16116);
   max_calc_reg_comparator_fourth_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx39793, D=>nx29241, CLK=>clk);
   ix29242 : oai21 port map ( Y=>nx29241, A0=>nx39793, A1=>nx41633, B0=>
      nx39796);
   ix39797 : nand03 port map ( Y=>nx39796, A0=>label_8_output_6, A1=>nx42643, 
      A2=>nx41633);
   ix29252 : oai21 port map ( Y=>nx29251, A0=>nx39800, A1=>nx41633, B0=>
      nx39802);
   max_calc_reg_comparator_fourth_inp1_6 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_6, QB=>nx39800, D=>nx29251, CLK=>clk);
   ix39803 : nand03 port map ( Y=>nx39802, A0=>label_7_output_6, A1=>nx42645, 
      A2=>nx41633);
   ix16117 : oai22 port map ( Y=>nx16116, A0=>nx39806, A1=>nx39819, B0=>
      max_calc_comparator_fourth_inp2_5, B1=>nx39814);
   ix29262 : oai21 port map ( Y=>nx29261, A0=>nx39810, A1=>nx41633, B0=>
      nx39812);
   max_calc_reg_comparator_fourth_inp2_5 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_5, QB=>nx39810, D=>nx29261, CLK=>clk);
   max_calc_reg_comparator_fourth_inp1_5 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_5, QB=>nx39814, D=>nx29271, CLK=>clk);
   ix29272 : oai21 port map ( Y=>nx29271, A0=>nx39814, A1=>nx41635, B0=>
      nx39817);
   ix39820 : aoi22 port map ( Y=>nx39819, A0=>nx39821, A1=>
      max_calc_comparator_fourth_inp1_4, B0=>nx15982, B1=>nx16100);
   max_calc_reg_comparator_fourth_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx39821, D=>nx29281, CLK=>clk);
   ix29282 : oai21 port map ( Y=>nx29281, A0=>nx39821, A1=>nx41635, B0=>
      nx39824);
   ix39825 : nand03 port map ( Y=>nx39824, A0=>label_8_output_4, A1=>nx42645, 
      A2=>nx41635);
   ix29292 : oai21 port map ( Y=>nx29291, A0=>nx39828, A1=>nx41635, B0=>
      nx39830);
   max_calc_reg_comparator_fourth_inp1_4 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_4, QB=>nx39828, D=>nx29291, CLK=>clk);
   ix39831 : nand03 port map ( Y=>nx39830, A0=>label_7_output_4, A1=>nx42645, 
      A2=>nx41635);
   ix16101 : oai22 port map ( Y=>nx16100, A0=>nx39834, A1=>nx39847, B0=>
      max_calc_comparator_fourth_inp2_3, B1=>nx39842);
   ix29302 : oai21 port map ( Y=>nx29301, A0=>nx39838, A1=>nx41637, B0=>
      nx39840);
   max_calc_reg_comparator_fourth_inp2_3 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_3, QB=>nx39838, D=>nx29301, CLK=>clk);
   max_calc_reg_comparator_fourth_inp1_3 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_3, QB=>nx39842, D=>nx29311, CLK=>clk);
   ix29312 : oai21 port map ( Y=>nx29311, A0=>nx39842, A1=>nx41637, B0=>
      nx39845);
   ix39848 : aoi22 port map ( Y=>nx39847, A0=>nx39849, A1=>
      max_calc_comparator_fourth_inp1_2, B0=>nx16026, B1=>nx16084);
   max_calc_reg_comparator_fourth_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx39849, D=>nx29321, CLK=>clk);
   ix29322 : oai21 port map ( Y=>nx29321, A0=>nx39849, A1=>nx41637, B0=>
      nx39852);
   ix39853 : nand03 port map ( Y=>nx39852, A0=>label_8_output_2, A1=>nx42647, 
      A2=>nx41637);
   ix29332 : oai21 port map ( Y=>nx29331, A0=>nx39856, A1=>nx41637, B0=>
      nx39858);
   max_calc_reg_comparator_fourth_inp1_2 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_2, QB=>nx39856, D=>nx29331, CLK=>clk);
   ix39859 : nand03 port map ( Y=>nx39858, A0=>label_7_output_2, A1=>nx42647, 
      A2=>nx41639);
   ix16085 : oai21 port map ( Y=>nx16084, A0=>
      max_calc_comparator_fourth_inp2_1, A1=>nx39868, B0=>nx39873);
   ix29342 : oai21 port map ( Y=>nx29341, A0=>nx39864, A1=>nx41639, B0=>
      nx39866);
   max_calc_reg_comparator_fourth_inp2_1 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_1, QB=>nx39864, D=>nx29341, CLK=>clk);
   max_calc_reg_comparator_fourth_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx39868, D=>nx29351, CLK=>clk);
   ix29352 : oai21 port map ( Y=>nx29351, A0=>nx39868, A1=>nx41639, B0=>
      nx39871);
   ix39874 : oai21 port map ( Y=>nx39873, A0=>nx39875, A1=>
      max_calc_comparator_fourth_inp1_0, B0=>nx16048);
   max_calc_reg_comparator_fourth_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx39875, D=>nx29361, CLK=>clk);
   ix29362 : oai21 port map ( Y=>nx29361, A0=>nx39875, A1=>nx41639, B0=>
      nx39878);
   ix39879 : nand03 port map ( Y=>nx39878, A0=>label_8_output_0, A1=>nx42647, 
      A2=>nx41639);
   ix29372 : oai21 port map ( Y=>nx29371, A0=>nx39882, A1=>nx41641, B0=>
      nx39884);
   max_calc_reg_comparator_fourth_inp1_0 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_0, QB=>nx39882, D=>nx29371, CLK=>clk);
   ix39885 : nand03 port map ( Y=>nx39884, A0=>label_7_output_0, A1=>nx42647, 
      A2=>nx41641);
   ix29402 : oai21 port map ( Y=>nx29401, A0=>nx39890, A1=>nx41641, B0=>
      nx39892);
   max_calc_reg_comparator_fourth_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx39890, D=>nx29401, CLK=>clk);
   lat_label_8_input_15 : latch port map ( Q=>label_8_input_15, D=>nx16210, 
      CLK=>nx41705);
   reg_label_8_input_state_machine_15 : dffr port map ( Q=>
      label_8_input_state_machine_15, QB=>OPEN, D=>nx29381, CLK=>clk, R=>rst
   );
   ix16207 : xnor2 port map ( Y=>nx16206, A0=>nx39902, A1=>nx16204);
   ix39903 : aoi22 port map ( Y=>nx39902, A0=>label_8_output_14, A1=>
      booth_booth_integration_output_7_26, B0=>nx15732, B1=>nx15734);
   labelsregfile_label8_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_8_output_15, QB=>nx39906, D=>nx29391, CLK=>clk, R=>rst);
   ix29432 : oai21 port map ( Y=>nx29431, A0=>nx39910, A1=>nx41641, B0=>
      nx39912);
   max_calc_reg_comparator_fourth_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx39910, D=>nx29431, CLK=>clk);
   lat_label_7_input_15 : latch port map ( Q=>label_7_input_15, D=>nx16252, 
      CLK=>nx41705);
   reg_label_7_input_state_machine_15 : dffr port map ( Q=>
      label_7_input_state_machine_15, QB=>OPEN, D=>nx29411, CLK=>clk, R=>rst
   );
   ix16249 : xnor2 port map ( Y=>nx16248, A0=>nx39922, A1=>nx16246);
   ix39923 : aoi22 port map ( Y=>nx39922, A0=>label_7_output_14, A1=>
      booth_booth_integration_output_6_26, B0=>nx14416, B1=>nx14418);
   labelsregfile_label7_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_7_output_15, QB=>nx39926, D=>nx29421, CLK=>clk, R=>rst);
   ix17605 : xnor2 port map ( Y=>nx17604, A0=>nx39930, A1=>nx17602);
   ix39931 : aoi22 port map ( Y=>nx39930, A0=>nx37785, A1=>
      max_calc_comparator_second_inp1_14, B0=>nx16310, B1=>nx17456);
   ix17457 : oai22 port map ( Y=>nx17456, A0=>nx39934, A1=>nx39957, B0=>
      max_calc_comparator_second_inp2_13, B1=>nx39947);
   ix29472 : oai21 port map ( Y=>nx29471, A0=>nx39938, A1=>nx41643, B0=>
      nx39940);
   max_calc_reg_comparator_second_inp2_13 : dff port map ( Q=>
      max_calc_comparator_second_inp2_13, QB=>nx39938, D=>nx29471, CLK=>clk
   );
   ix39941 : nand03 port map ( Y=>nx39940, A0=>nx42819, A1=>nx16336, A2=>
      nx41643);
   max_calc_reg_ans4_13 : dff port map ( Q=>max_calc_ans4_13, QB=>OPEN, D=>
      nx29461, CLK=>clk);
   ix29462 : ao32 port map ( Y=>nx29461, A0=>nx42229, A1=>nx16322, A2=>
      nx41811, B0=>max_calc_ans4_13, B1=>nx42679);
   max_calc_reg_comparator_second_inp1_13 : dff port map ( Q=>
      max_calc_comparator_second_inp1_13, QB=>nx39947, D=>nx29491, CLK=>clk
   );
   ix29492 : oai21 port map ( Y=>nx29491, A0=>nx39947, A1=>nx41643, B0=>
      nx39950);
   ix39951 : nand03 port map ( Y=>nx39950, A0=>nx42229, A1=>nx16372, A2=>
      nx41643);
   max_calc_reg_ans3_13 : dff port map ( Q=>max_calc_ans3_13, QB=>OPEN, D=>
      nx29481, CLK=>clk);
   ix29482 : ao32 port map ( Y=>nx29481, A0=>nx42229, A1=>nx16358, A2=>
      nx41811, B0=>max_calc_ans3_13, B1=>nx42679);
   ix39958 : aoi22 port map ( Y=>nx39957, A0=>nx39959, A1=>
      max_calc_comparator_second_inp1_12, B0=>nx16458, B1=>nx17440);
   max_calc_reg_comparator_second_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx39959, D=>nx29511, CLK=>clk);
   ix29512 : oai21 port map ( Y=>nx29511, A0=>nx39959, A1=>nx41643, B0=>
      nx39962);
   ix39963 : nand03 port map ( Y=>nx39962, A0=>nx42229, A1=>nx16410, A2=>
      nx41643);
   max_calc_reg_ans4_12 : dff port map ( Q=>max_calc_ans4_12, QB=>OPEN, D=>
      nx29501, CLK=>clk);
   ix29502 : ao32 port map ( Y=>nx29501, A0=>nx42229, A1=>nx16396, A2=>
      nx41813, B0=>max_calc_ans4_12, B1=>nx42679);
   ix29532 : oai21 port map ( Y=>nx29531, A0=>nx39971, A1=>nx41643, B0=>
      nx39973);
   max_calc_reg_comparator_second_inp1_12 : dff port map ( Q=>
      max_calc_comparator_second_inp1_12, QB=>nx39971, D=>nx29531, CLK=>clk
   );
   ix39974 : nand03 port map ( Y=>nx39973, A0=>nx42229, A1=>nx16446, A2=>
      nx41645);
   max_calc_reg_ans3_12 : dff port map ( Q=>max_calc_ans3_12, QB=>OPEN, D=>
      nx29521, CLK=>clk);
   ix29522 : ao32 port map ( Y=>nx29521, A0=>nx42229, A1=>nx16432, A2=>
      nx41813, B0=>max_calc_ans3_12, B1=>nx42679);
   ix17441 : oai22 port map ( Y=>nx17440, A0=>nx39982, A1=>nx40005, B0=>
      max_calc_comparator_second_inp2_11, B1=>nx39995);
   ix29552 : oai21 port map ( Y=>nx29551, A0=>nx39986, A1=>nx41645, B0=>
      nx39988);
   max_calc_reg_comparator_second_inp2_11 : dff port map ( Q=>
      max_calc_comparator_second_inp2_11, QB=>nx39986, D=>nx29551, CLK=>clk
   );
   ix39989 : nand03 port map ( Y=>nx39988, A0=>nx42231, A1=>nx16484, A2=>
      nx41645);
   max_calc_reg_ans4_11 : dff port map ( Q=>max_calc_ans4_11, QB=>OPEN, D=>
      nx29541, CLK=>clk);
   ix29542 : ao32 port map ( Y=>nx29541, A0=>nx42231, A1=>nx16470, A2=>
      nx41813, B0=>max_calc_ans4_11, B1=>nx42679);
   max_calc_reg_comparator_second_inp1_11 : dff port map ( Q=>
      max_calc_comparator_second_inp1_11, QB=>nx39995, D=>nx29571, CLK=>clk
   );
   ix29572 : oai21 port map ( Y=>nx29571, A0=>nx39995, A1=>nx41645, B0=>
      nx39998);
   ix39999 : nand03 port map ( Y=>nx39998, A0=>nx42231, A1=>nx16520, A2=>
      nx41645);
   max_calc_reg_ans3_11 : dff port map ( Q=>max_calc_ans3_11, QB=>OPEN, D=>
      nx29561, CLK=>clk);
   ix29562 : ao32 port map ( Y=>nx29561, A0=>nx42231, A1=>nx16506, A2=>
      nx41813, B0=>max_calc_ans3_11, B1=>nx42681);
   ix40006 : aoi22 port map ( Y=>nx40005, A0=>nx40007, A1=>
      max_calc_comparator_second_inp1_10, B0=>nx16606, B1=>nx17424);
   max_calc_reg_comparator_second_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx40007, D=>nx29591, CLK=>clk);
   ix29592 : oai21 port map ( Y=>nx29591, A0=>nx40007, A1=>nx41645, B0=>
      nx40010);
   ix40011 : nand03 port map ( Y=>nx40010, A0=>nx42231, A1=>nx16558, A2=>
      nx41645);
   max_calc_reg_ans4_10 : dff port map ( Q=>max_calc_ans4_10, QB=>OPEN, D=>
      nx29581, CLK=>clk);
   ix29582 : ao32 port map ( Y=>nx29581, A0=>nx42231, A1=>nx16544, A2=>
      nx41813, B0=>max_calc_ans4_10, B1=>nx42681);
   ix29612 : oai21 port map ( Y=>nx29611, A0=>nx40019, A1=>nx41647, B0=>
      nx40021);
   max_calc_reg_comparator_second_inp1_10 : dff port map ( Q=>
      max_calc_comparator_second_inp1_10, QB=>nx40019, D=>nx29611, CLK=>clk
   );
   ix40022 : nand03 port map ( Y=>nx40021, A0=>nx42231, A1=>nx16594, A2=>
      nx41647);
   max_calc_reg_ans3_10 : dff port map ( Q=>max_calc_ans3_10, QB=>OPEN, D=>
      nx29601, CLK=>clk);
   ix29602 : ao32 port map ( Y=>nx29601, A0=>nx42233, A1=>nx16580, A2=>
      nx41813, B0=>max_calc_ans3_10, B1=>nx42681);
   ix17425 : oai22 port map ( Y=>nx17424, A0=>nx40030, A1=>nx40053, B0=>
      max_calc_comparator_second_inp2_9, B1=>nx40043);
   ix29632 : oai21 port map ( Y=>nx29631, A0=>nx40034, A1=>nx41647, B0=>
      nx40036);
   max_calc_reg_comparator_second_inp2_9 : dff port map ( Q=>
      max_calc_comparator_second_inp2_9, QB=>nx40034, D=>nx29631, CLK=>clk);
   ix40037 : nand03 port map ( Y=>nx40036, A0=>nx42233, A1=>nx16632, A2=>
      nx41647);
   max_calc_reg_ans4_9 : dff port map ( Q=>max_calc_ans4_9, QB=>OPEN, D=>
      nx29621, CLK=>clk);
   ix29622 : ao32 port map ( Y=>nx29621, A0=>nx42233, A1=>nx16618, A2=>
      nx41813, B0=>max_calc_ans4_9, B1=>nx42681);
   max_calc_reg_comparator_second_inp1_9 : dff port map ( Q=>
      max_calc_comparator_second_inp1_9, QB=>nx40043, D=>nx29651, CLK=>clk);
   ix29652 : oai21 port map ( Y=>nx29651, A0=>nx40043, A1=>nx41647, B0=>
      nx40046);
   ix40047 : nand03 port map ( Y=>nx40046, A0=>nx42233, A1=>nx16668, A2=>
      nx41647);
   max_calc_reg_ans3_9 : dff port map ( Q=>max_calc_ans3_9, QB=>OPEN, D=>
      nx29641, CLK=>clk);
   ix29642 : ao32 port map ( Y=>nx29641, A0=>nx42233, A1=>nx16654, A2=>
      nx41815, B0=>max_calc_ans3_9, B1=>nx42681);
   ix40054 : aoi22 port map ( Y=>nx40053, A0=>nx40055, A1=>
      max_calc_comparator_second_inp1_8, B0=>nx16754, B1=>nx17408);
   max_calc_reg_comparator_second_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx40055, D=>nx29671, CLK=>clk);
   ix29672 : oai21 port map ( Y=>nx29671, A0=>nx40055, A1=>nx41647, B0=>
      nx40058);
   ix40059 : nand03 port map ( Y=>nx40058, A0=>nx42233, A1=>nx16706, A2=>
      nx41649);
   max_calc_reg_ans4_8 : dff port map ( Q=>max_calc_ans4_8, QB=>OPEN, D=>
      nx29661, CLK=>clk);
   ix29662 : ao32 port map ( Y=>nx29661, A0=>nx42233, A1=>nx16692, A2=>
      nx41815, B0=>max_calc_ans4_8, B1=>nx42681);
   ix29692 : oai21 port map ( Y=>nx29691, A0=>nx40067, A1=>nx41649, B0=>
      nx40069);
   max_calc_reg_comparator_second_inp1_8 : dff port map ( Q=>
      max_calc_comparator_second_inp1_8, QB=>nx40067, D=>nx29691, CLK=>clk);
   ix40070 : nand03 port map ( Y=>nx40069, A0=>nx42235, A1=>nx16742, A2=>
      nx41649);
   max_calc_reg_ans3_8 : dff port map ( Q=>max_calc_ans3_8, QB=>OPEN, D=>
      nx29681, CLK=>clk);
   ix29682 : ao32 port map ( Y=>nx29681, A0=>nx42235, A1=>nx16728, A2=>
      nx41815, B0=>max_calc_ans3_8, B1=>nx42681);
   ix17409 : oai22 port map ( Y=>nx17408, A0=>nx40078, A1=>nx40101, B0=>
      max_calc_comparator_second_inp2_7, B1=>nx40091);
   ix29712 : oai21 port map ( Y=>nx29711, A0=>nx40082, A1=>nx41649, B0=>
      nx40084);
   max_calc_reg_comparator_second_inp2_7 : dff port map ( Q=>
      max_calc_comparator_second_inp2_7, QB=>nx40082, D=>nx29711, CLK=>clk);
   ix40085 : nand03 port map ( Y=>nx40084, A0=>nx42235, A1=>nx16780, A2=>
      nx41649);
   max_calc_reg_ans4_7 : dff port map ( Q=>max_calc_ans4_7, QB=>OPEN, D=>
      nx29701, CLK=>clk);
   ix29702 : ao32 port map ( Y=>nx29701, A0=>nx42235, A1=>nx16766, A2=>
      nx41815, B0=>max_calc_ans4_7, B1=>nx42683);
   max_calc_reg_comparator_second_inp1_7 : dff port map ( Q=>
      max_calc_comparator_second_inp1_7, QB=>nx40091, D=>nx29731, CLK=>clk);
   ix29732 : oai21 port map ( Y=>nx29731, A0=>nx40091, A1=>nx41649, B0=>
      nx40094);
   ix40095 : nand03 port map ( Y=>nx40094, A0=>nx42235, A1=>nx16816, A2=>
      nx41649);
   max_calc_reg_ans3_7 : dff port map ( Q=>max_calc_ans3_7, QB=>OPEN, D=>
      nx29721, CLK=>clk);
   ix29722 : ao32 port map ( Y=>nx29721, A0=>nx42235, A1=>nx16802, A2=>
      nx41815, B0=>max_calc_ans3_7, B1=>nx42683);
   ix40102 : aoi22 port map ( Y=>nx40101, A0=>nx40103, A1=>
      max_calc_comparator_second_inp1_6, B0=>nx16902, B1=>nx17392);
   max_calc_reg_comparator_second_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx40103, D=>nx29751, CLK=>clk);
   ix29752 : oai21 port map ( Y=>nx29751, A0=>nx40103, A1=>nx41651, B0=>
      nx40106);
   ix40107 : nand03 port map ( Y=>nx40106, A0=>nx42235, A1=>nx16854, A2=>
      nx41651);
   max_calc_reg_ans4_6 : dff port map ( Q=>max_calc_ans4_6, QB=>OPEN, D=>
      nx29741, CLK=>clk);
   ix29742 : ao32 port map ( Y=>nx29741, A0=>nx42237, A1=>nx16840, A2=>
      nx41815, B0=>max_calc_ans4_6, B1=>nx42683);
   ix29772 : oai21 port map ( Y=>nx29771, A0=>nx40115, A1=>nx41651, B0=>
      nx40117);
   max_calc_reg_comparator_second_inp1_6 : dff port map ( Q=>
      max_calc_comparator_second_inp1_6, QB=>nx40115, D=>nx29771, CLK=>clk);
   ix40118 : nand03 port map ( Y=>nx40117, A0=>nx42237, A1=>nx16890, A2=>
      nx41651);
   max_calc_reg_ans3_6 : dff port map ( Q=>max_calc_ans3_6, QB=>OPEN, D=>
      nx29761, CLK=>clk);
   ix29762 : ao32 port map ( Y=>nx29761, A0=>nx42237, A1=>nx16876, A2=>
      nx41815, B0=>max_calc_ans3_6, B1=>nx42683);
   ix17393 : oai22 port map ( Y=>nx17392, A0=>nx40126, A1=>nx40149, B0=>
      max_calc_comparator_second_inp2_5, B1=>nx40139);
   ix29792 : oai21 port map ( Y=>nx29791, A0=>nx40130, A1=>nx41651, B0=>
      nx40132);
   max_calc_reg_comparator_second_inp2_5 : dff port map ( Q=>
      max_calc_comparator_second_inp2_5, QB=>nx40130, D=>nx29791, CLK=>clk);
   ix40133 : nand03 port map ( Y=>nx40132, A0=>nx42237, A1=>nx16928, A2=>
      nx41651);
   max_calc_reg_ans4_5 : dff port map ( Q=>max_calc_ans4_5, QB=>OPEN, D=>
      nx29781, CLK=>clk);
   ix29782 : ao32 port map ( Y=>nx29781, A0=>nx42237, A1=>nx16914, A2=>
      nx41817, B0=>max_calc_ans4_5, B1=>nx42683);
   max_calc_reg_comparator_second_inp1_5 : dff port map ( Q=>
      max_calc_comparator_second_inp1_5, QB=>nx40139, D=>nx29811, CLK=>clk);
   ix29812 : oai21 port map ( Y=>nx29811, A0=>nx40139, A1=>nx41651, B0=>
      nx40142);
   ix40143 : nand03 port map ( Y=>nx40142, A0=>nx42237, A1=>nx16964, A2=>
      nx41653);
   max_calc_reg_ans3_5 : dff port map ( Q=>max_calc_ans3_5, QB=>OPEN, D=>
      nx29801, CLK=>clk);
   ix29802 : ao32 port map ( Y=>nx29801, A0=>nx42237, A1=>nx16950, A2=>
      nx41817, B0=>max_calc_ans3_5, B1=>nx42683);
   ix40150 : aoi22 port map ( Y=>nx40149, A0=>nx40151, A1=>
      max_calc_comparator_second_inp1_4, B0=>nx17050, B1=>nx17376);
   max_calc_reg_comparator_second_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx40151, D=>nx29831, CLK=>clk);
   ix29832 : oai21 port map ( Y=>nx29831, A0=>nx40151, A1=>nx41653, B0=>
      nx40154);
   ix40155 : nand03 port map ( Y=>nx40154, A0=>nx42239, A1=>nx17002, A2=>
      nx41653);
   max_calc_reg_ans4_4 : dff port map ( Q=>max_calc_ans4_4, QB=>OPEN, D=>
      nx29821, CLK=>clk);
   ix29822 : ao32 port map ( Y=>nx29821, A0=>nx42239, A1=>nx16988, A2=>
      nx41817, B0=>max_calc_ans4_4, B1=>nx42683);
   ix29852 : oai21 port map ( Y=>nx29851, A0=>nx40163, A1=>nx41653, B0=>
      nx40165);
   max_calc_reg_comparator_second_inp1_4 : dff port map ( Q=>
      max_calc_comparator_second_inp1_4, QB=>nx40163, D=>nx29851, CLK=>clk);
   ix40166 : nand03 port map ( Y=>nx40165, A0=>nx42239, A1=>nx17038, A2=>
      nx41653);
   max_calc_reg_ans3_4 : dff port map ( Q=>max_calc_ans3_4, QB=>OPEN, D=>
      nx29841, CLK=>clk);
   ix29842 : ao32 port map ( Y=>nx29841, A0=>nx42239, A1=>nx17024, A2=>
      nx41817, B0=>max_calc_ans3_4, B1=>nx42685);
   ix17377 : oai22 port map ( Y=>nx17376, A0=>nx40174, A1=>nx40197, B0=>
      max_calc_comparator_second_inp2_3, B1=>nx40187);
   ix29872 : oai21 port map ( Y=>nx29871, A0=>nx40178, A1=>nx41653, B0=>
      nx40180);
   max_calc_reg_comparator_second_inp2_3 : dff port map ( Q=>
      max_calc_comparator_second_inp2_3, QB=>nx40178, D=>nx29871, CLK=>clk);
   ix40181 : nand03 port map ( Y=>nx40180, A0=>nx42239, A1=>nx17076, A2=>
      nx41653);
   max_calc_reg_ans4_3 : dff port map ( Q=>max_calc_ans4_3, QB=>OPEN, D=>
      nx29861, CLK=>clk);
   ix29862 : ao32 port map ( Y=>nx29861, A0=>nx42239, A1=>nx17062, A2=>
      nx41817, B0=>max_calc_ans4_3, B1=>nx42685);
   max_calc_reg_comparator_second_inp1_3 : dff port map ( Q=>
      max_calc_comparator_second_inp1_3, QB=>nx40187, D=>nx29891, CLK=>clk);
   ix29892 : oai21 port map ( Y=>nx29891, A0=>nx40187, A1=>nx41655, B0=>
      nx40190);
   ix40191 : nand03 port map ( Y=>nx40190, A0=>nx42239, A1=>nx17112, A2=>
      nx41655);
   max_calc_reg_ans3_3 : dff port map ( Q=>max_calc_ans3_3, QB=>OPEN, D=>
      nx29881, CLK=>clk);
   ix29882 : ao32 port map ( Y=>nx29881, A0=>nx42241, A1=>nx17098, A2=>
      nx41817, B0=>max_calc_ans3_3, B1=>nx42685);
   ix40198 : aoi22 port map ( Y=>nx40197, A0=>nx40199, A1=>
      max_calc_comparator_second_inp1_2, B0=>nx17198, B1=>nx17360);
   max_calc_reg_comparator_second_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx40199, D=>nx29911, CLK=>clk);
   ix29912 : oai21 port map ( Y=>nx29911, A0=>nx40199, A1=>nx41655, B0=>
      nx40202);
   ix40203 : nand03 port map ( Y=>nx40202, A0=>nx42241, A1=>nx17150, A2=>
      nx41655);
   max_calc_reg_ans4_2 : dff port map ( Q=>max_calc_ans4_2, QB=>OPEN, D=>
      nx29901, CLK=>clk);
   ix29902 : ao32 port map ( Y=>nx29901, A0=>nx42241, A1=>nx17136, A2=>
      nx41817, B0=>max_calc_ans4_2, B1=>nx42685);
   ix29932 : oai21 port map ( Y=>nx29931, A0=>nx40211, A1=>nx41655, B0=>
      nx40213);
   max_calc_reg_comparator_second_inp1_2 : dff port map ( Q=>
      max_calc_comparator_second_inp1_2, QB=>nx40211, D=>nx29931, CLK=>clk);
   ix40214 : nand03 port map ( Y=>nx40213, A0=>nx42241, A1=>nx17186, A2=>
      nx41655);
   max_calc_reg_ans3_2 : dff port map ( Q=>max_calc_ans3_2, QB=>OPEN, D=>
      nx29921, CLK=>clk);
   ix29922 : ao32 port map ( Y=>nx29921, A0=>nx42241, A1=>nx17172, A2=>
      nx41819, B0=>max_calc_ans3_2, B1=>nx42685);
   ix17361 : oai21 port map ( Y=>nx17360, A0=>
      max_calc_comparator_second_inp2_1, A1=>nx40233, B0=>nx40243);
   ix29952 : oai21 port map ( Y=>nx29951, A0=>nx40224, A1=>nx41655, B0=>
      nx40226);
   max_calc_reg_comparator_second_inp2_1 : dff port map ( Q=>
      max_calc_comparator_second_inp2_1, QB=>nx40224, D=>nx29951, CLK=>clk);
   ix40227 : nand03 port map ( Y=>nx40226, A0=>nx42241, A1=>nx17224, A2=>
      nx41657);
   max_calc_reg_ans4_1 : dff port map ( Q=>max_calc_ans4_1, QB=>OPEN, D=>
      nx29941, CLK=>clk);
   ix29942 : ao32 port map ( Y=>nx29941, A0=>nx42241, A1=>nx17210, A2=>
      nx41819, B0=>max_calc_ans4_1, B1=>nx42685);
   max_calc_reg_comparator_second_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx40233, D=>nx29971, CLK=>clk);
   ix29972 : oai21 port map ( Y=>nx29971, A0=>nx40233, A1=>nx41657, B0=>
      nx40236);
   ix40237 : nand03 port map ( Y=>nx40236, A0=>nx42243, A1=>nx17260, A2=>
      nx41657);
   max_calc_reg_ans3_1 : dff port map ( Q=>max_calc_ans3_1, QB=>OPEN, D=>
      nx29961, CLK=>clk);
   ix29962 : ao32 port map ( Y=>nx29961, A0=>nx42243, A1=>nx17246, A2=>
      nx41819, B0=>max_calc_ans3_1, B1=>nx42685);
   ix40244 : oai21 port map ( Y=>nx40243, A0=>nx40245, A1=>
      max_calc_comparator_second_inp1_0, B0=>nx17272);
   max_calc_reg_comparator_second_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx40245, D=>nx29991, CLK=>clk);
   ix29992 : oai21 port map ( Y=>nx29991, A0=>nx40245, A1=>nx41657, B0=>
      nx40248);
   ix40249 : nand03 port map ( Y=>nx40248, A0=>nx42243, A1=>nx17298, A2=>
      nx41657);
   max_calc_reg_ans4_0 : dff port map ( Q=>max_calc_ans4_0, QB=>OPEN, D=>
      nx29981, CLK=>clk);
   ix29982 : ao32 port map ( Y=>nx29981, A0=>nx42243, A1=>nx17284, A2=>
      nx41819, B0=>max_calc_ans4_0, B1=>nx42687);
   ix30012 : oai21 port map ( Y=>nx30011, A0=>nx40257, A1=>nx41657, B0=>
      nx40259);
   max_calc_reg_comparator_second_inp1_0 : dff port map ( Q=>
      max_calc_comparator_second_inp1_0, QB=>nx40257, D=>nx30011, CLK=>clk);
   ix40260 : nand03 port map ( Y=>nx40259, A0=>nx42243, A1=>nx17334, A2=>
      nx41657);
   max_calc_reg_ans3_0 : dff port map ( Q=>max_calc_ans3_0, QB=>OPEN, D=>
      nx30001, CLK=>clk);
   ix30002 : ao32 port map ( Y=>nx30001, A0=>nx42243, A1=>nx17320, A2=>
      nx41819, B0=>max_calc_ans3_0, B1=>nx42687);
   ix30052 : oai21 port map ( Y=>nx30051, A0=>nx40270, A1=>nx41659, B0=>
      nx40272);
   max_calc_reg_comparator_second_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx40270, D=>nx30051, CLK=>clk);
   ix40273 : nand03 port map ( Y=>nx40272, A0=>nx42243, A1=>nx17522, A2=>
      nx41659);
   lat_label_4_input_15 : latch port map ( Q=>label_4_input_15, D=>nx17486, 
      CLK=>nx41705);
   reg_label_4_input_state_machine_15 : dffr port map ( Q=>
      label_4_input_state_machine_15, QB=>OPEN, D=>nx30021, CLK=>clk, R=>rst
   );
   ix17483 : xnor2 port map ( Y=>nx17482, A0=>nx40283, A1=>nx17480);
   ix40284 : aoi22 port map ( Y=>nx40283, A0=>label_4_output_14, A1=>
      booth_booth_integration_output_3_26, B0=>nx13106, B1=>nx13108);
   labelsregfile_label4_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_4_output_15, QB=>nx40287, D=>nx30031, CLK=>clk, R=>rst);
   max_calc_reg_ans4_15 : dff port map ( Q=>max_calc_ans4_15, QB=>OPEN, D=>
      nx30041, CLK=>clk);
   ix30042 : ao32 port map ( Y=>nx30041, A0=>nx42245, A1=>nx17508, A2=>
      nx41819, B0=>max_calc_ans4_15, B1=>nx42687);
   ix30092 : oai21 port map ( Y=>nx30091, A0=>nx40295, A1=>nx41659, B0=>
      nx40297);
   max_calc_reg_comparator_second_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx40295, D=>nx30091, CLK=>clk);
   ix40298 : nand03 port map ( Y=>nx40297, A0=>nx42245, A1=>nx17590, A2=>
      nx41659);
   lat_label_3_input_15 : latch port map ( Q=>label_3_input_15, D=>nx17554, 
      CLK=>nx41705);
   reg_label_3_input_state_machine_15 : dffr port map ( Q=>
      label_3_input_state_machine_15, QB=>OPEN, D=>nx30061, CLK=>clk, R=>rst
   );
   ix17551 : xnor2 port map ( Y=>nx17550, A0=>nx40308, A1=>nx17548);
   ix40309 : aoi22 port map ( Y=>nx40308, A0=>label_3_output_14, A1=>
      booth_booth_integration_output_2_26, B0=>nx8604, B1=>nx8606);
   labelsregfile_label3_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_3_output_15, QB=>nx40312, D=>nx30071, CLK=>clk, R=>rst);
   max_calc_reg_ans3_15 : dff port map ( Q=>max_calc_ans3_15, QB=>OPEN, D=>
      nx30081, CLK=>clk);
   ix30082 : ao32 port map ( Y=>nx30081, A0=>nx42245, A1=>nx17576, A2=>
      nx41819, B0=>max_calc_ans3_15, B1=>nx42687);
   max_calc_reg_ans7_14 : dff port map ( Q=>max_calc_ans7_14, QB=>OPEN, D=>
      nx30441, CLK=>clk);
   max_calc_reg_ans8_14 : dff port map ( Q=>max_calc_ans8_14, QB=>OPEN, D=>
      nx30431, CLK=>clk);
   ix20115 : xnor2 port map ( Y=>nx18605, A0=>nx40328, A1=>nx20112);
   ix40329 : aoi22 port map ( Y=>nx40328, A0=>nx40326, A1=>
      max_calc_comparator_first_inp1_14, B0=>nx18164, B1=>nx19918);
   ix19919 : oai22 port map ( Y=>nx19918, A0=>nx40332, A1=>nx40367, B0=>
      max_calc_comparator_first_inp2_13, B1=>nx40364);
   max_calc_reg_comparator_first_inp2_13 : dff port map ( Q=>
      max_calc_comparator_first_inp2_13, QB=>OPEN, D=>nx30531, CLK=>clk);
   max_calc_reg_ans2_13 : dff port map ( Q=>max_calc_ans2_13, QB=>OPEN, D=>
      nx30461, CLK=>clk);
   max_calc_reg_ans7_13 : dff port map ( Q=>max_calc_ans7_13, QB=>OPEN, D=>
      nx30521, CLK=>clk);
   max_calc_reg_ans8_13 : dff port map ( Q=>max_calc_ans8_13, QB=>OPEN, D=>
      nx30511, CLK=>clk);
   max_calc_reg_comparator_first_inp1_13 : dff port map ( Q=>
      max_calc_comparator_first_inp1_13, QB=>nx40364, D=>nx30501, CLK=>clk);
   max_calc_reg_ans1_13 : dff port map ( Q=>max_calc_ans1_13, QB=>OPEN, D=>
      nx30471, CLK=>clk);
   max_calc_reg_ans6_13 : dff port map ( Q=>max_calc_ans6_13, QB=>OPEN, D=>
      nx30481, CLK=>clk);
   max_calc_reg_ans5_13 : dff port map ( Q=>max_calc_ans5_13, QB=>OPEN, D=>
      nx30491, CLK=>clk);
   ix40368 : aoi22 port map ( Y=>nx40367, A0=>nx40369, A1=>
      max_calc_comparator_first_inp1_12, B0=>nx18408, B1=>nx19902);
   max_calc_reg_ans2_12 : dff port map ( Q=>max_calc_ans2_12, QB=>OPEN, D=>
      nx30541, CLK=>clk);
   max_calc_reg_ans7_12 : dff port map ( Q=>max_calc_ans7_12, QB=>OPEN, D=>
      nx30601, CLK=>clk);
   max_calc_reg_ans8_12 : dff port map ( Q=>max_calc_ans8_12, QB=>OPEN, D=>
      nx30591, CLK=>clk);
   max_calc_reg_comparator_first_inp1_12 : dff port map ( Q=>
      max_calc_comparator_first_inp1_12, QB=>OPEN, D=>nx30581, CLK=>clk);
   max_calc_reg_ans1_12 : dff port map ( Q=>max_calc_ans1_12, QB=>OPEN, D=>
      nx30551, CLK=>clk);
   max_calc_reg_ans6_12 : dff port map ( Q=>max_calc_ans6_12, QB=>OPEN, D=>
      nx30561, CLK=>clk);
   max_calc_reg_ans5_12 : dff port map ( Q=>max_calc_ans5_12, QB=>OPEN, D=>
      nx30571, CLK=>clk);
   max_calc_reg_comparator_first_inp2_12 : dff port map ( Q=>
      max_calc_comparator_first_inp2_12, QB=>nx40369, D=>nx30611, CLK=>clk);
   ix19903 : oai22 port map ( Y=>nx19902, A0=>nx40405, A1=>nx40440, B0=>
      max_calc_comparator_first_inp2_11, B1=>nx40437);
   max_calc_reg_comparator_first_inp2_11 : dff port map ( Q=>
      max_calc_comparator_first_inp2_11, QB=>OPEN, D=>nx30691, CLK=>clk);
   max_calc_reg_ans2_11 : dff port map ( Q=>max_calc_ans2_11, QB=>OPEN, D=>
      nx30621, CLK=>clk);
   max_calc_reg_ans7_11 : dff port map ( Q=>max_calc_ans7_11, QB=>OPEN, D=>
      nx30681, CLK=>clk);
   max_calc_reg_ans8_11 : dff port map ( Q=>max_calc_ans8_11, QB=>OPEN, D=>
      nx30671, CLK=>clk);
   max_calc_reg_comparator_first_inp1_11 : dff port map ( Q=>
      max_calc_comparator_first_inp1_11, QB=>nx40437, D=>nx30661, CLK=>clk);
   max_calc_reg_ans1_11 : dff port map ( Q=>max_calc_ans1_11, QB=>OPEN, D=>
      nx30631, CLK=>clk);
   max_calc_reg_ans6_11 : dff port map ( Q=>max_calc_ans6_11, QB=>OPEN, D=>
      nx30641, CLK=>clk);
   max_calc_reg_ans5_11 : dff port map ( Q=>max_calc_ans5_11, QB=>OPEN, D=>
      nx30651, CLK=>clk);
   ix40441 : aoi22 port map ( Y=>nx40440, A0=>nx40442, A1=>
      max_calc_comparator_first_inp1_10, B0=>nx18652, B1=>nx19886);
   max_calc_reg_ans2_10 : dff port map ( Q=>max_calc_ans2_10, QB=>OPEN, D=>
      nx30701, CLK=>clk);
   max_calc_reg_ans7_10 : dff port map ( Q=>max_calc_ans7_10, QB=>OPEN, D=>
      nx30761, CLK=>clk);
   max_calc_reg_ans8_10 : dff port map ( Q=>max_calc_ans8_10, QB=>OPEN, D=>
      nx30751, CLK=>clk);
   max_calc_reg_comparator_first_inp1_10 : dff port map ( Q=>
      max_calc_comparator_first_inp1_10, QB=>OPEN, D=>nx30741, CLK=>clk);
   max_calc_reg_ans1_10 : dff port map ( Q=>max_calc_ans1_10, QB=>OPEN, D=>
      nx30711, CLK=>clk);
   max_calc_reg_ans6_10 : dff port map ( Q=>max_calc_ans6_10, QB=>OPEN, D=>
      nx30721, CLK=>clk);
   max_calc_reg_ans5_10 : dff port map ( Q=>max_calc_ans5_10, QB=>OPEN, D=>
      nx30731, CLK=>clk);
   max_calc_reg_comparator_first_inp2_10 : dff port map ( Q=>
      max_calc_comparator_first_inp2_10, QB=>nx40442, D=>nx30771, CLK=>clk);
   ix19887 : oai22 port map ( Y=>nx19886, A0=>nx40478, A1=>nx40513, B0=>
      max_calc_comparator_first_inp2_9, B1=>nx40510);
   max_calc_reg_comparator_first_inp2_9 : dff port map ( Q=>
      max_calc_comparator_first_inp2_9, QB=>OPEN, D=>nx30851, CLK=>clk);
   max_calc_reg_ans2_9 : dff port map ( Q=>max_calc_ans2_9, QB=>OPEN, D=>
      nx30781, CLK=>clk);
   max_calc_reg_ans7_9 : dff port map ( Q=>max_calc_ans7_9, QB=>OPEN, D=>
      nx30841, CLK=>clk);
   max_calc_reg_ans8_9 : dff port map ( Q=>max_calc_ans8_9, QB=>OPEN, D=>
      nx30831, CLK=>clk);
   max_calc_reg_comparator_first_inp1_9 : dff port map ( Q=>
      max_calc_comparator_first_inp1_9, QB=>nx40510, D=>nx30821, CLK=>clk);
   max_calc_reg_ans1_9 : dff port map ( Q=>max_calc_ans1_9, QB=>OPEN, D=>
      nx30791, CLK=>clk);
   max_calc_reg_ans6_9 : dff port map ( Q=>max_calc_ans6_9, QB=>OPEN, D=>
      nx30801, CLK=>clk);
   max_calc_reg_ans5_9 : dff port map ( Q=>max_calc_ans5_9, QB=>OPEN, D=>
      nx30811, CLK=>clk);
   ix40514 : aoi22 port map ( Y=>nx40513, A0=>nx40515, A1=>
      max_calc_comparator_first_inp1_8, B0=>nx18896, B1=>nx19870);
   max_calc_reg_ans2_8 : dff port map ( Q=>max_calc_ans2_8, QB=>OPEN, D=>
      nx30861, CLK=>clk);
   max_calc_reg_ans7_8 : dff port map ( Q=>max_calc_ans7_8, QB=>OPEN, D=>
      nx30921, CLK=>clk);
   max_calc_reg_ans8_8 : dff port map ( Q=>max_calc_ans8_8, QB=>OPEN, D=>
      nx30911, CLK=>clk);
   max_calc_reg_comparator_first_inp1_8 : dff port map ( Q=>
      max_calc_comparator_first_inp1_8, QB=>OPEN, D=>nx30901, CLK=>clk);
   max_calc_reg_ans1_8 : dff port map ( Q=>max_calc_ans1_8, QB=>OPEN, D=>
      nx30871, CLK=>clk);
   max_calc_reg_ans6_8 : dff port map ( Q=>max_calc_ans6_8, QB=>OPEN, D=>
      nx30881, CLK=>clk);
   max_calc_reg_ans5_8 : dff port map ( Q=>max_calc_ans5_8, QB=>OPEN, D=>
      nx30891, CLK=>clk);
   max_calc_reg_comparator_first_inp2_8 : dff port map ( Q=>
      max_calc_comparator_first_inp2_8, QB=>nx40515, D=>nx30931, CLK=>clk);
   ix19871 : oai22 port map ( Y=>nx19870, A0=>nx40551, A1=>nx40586, B0=>
      max_calc_comparator_first_inp2_7, B1=>nx40583);
   max_calc_reg_comparator_first_inp2_7 : dff port map ( Q=>
      max_calc_comparator_first_inp2_7, QB=>OPEN, D=>nx31011, CLK=>clk);
   max_calc_reg_ans2_7 : dff port map ( Q=>max_calc_ans2_7, QB=>OPEN, D=>
      nx30941, CLK=>clk);
   max_calc_reg_ans7_7 : dff port map ( Q=>max_calc_ans7_7, QB=>OPEN, D=>
      nx31001, CLK=>clk);
   max_calc_reg_ans8_7 : dff port map ( Q=>max_calc_ans8_7, QB=>OPEN, D=>
      nx30991, CLK=>clk);
   max_calc_reg_comparator_first_inp1_7 : dff port map ( Q=>
      max_calc_comparator_first_inp1_7, QB=>nx40583, D=>nx30981, CLK=>clk);
   max_calc_reg_ans1_7 : dff port map ( Q=>max_calc_ans1_7, QB=>OPEN, D=>
      nx30951, CLK=>clk);
   max_calc_reg_ans6_7 : dff port map ( Q=>max_calc_ans6_7, QB=>OPEN, D=>
      nx30961, CLK=>clk);
   max_calc_reg_ans5_7 : dff port map ( Q=>max_calc_ans5_7, QB=>OPEN, D=>
      nx30971, CLK=>clk);
   ix40587 : aoi22 port map ( Y=>nx40586, A0=>nx40588, A1=>
      max_calc_comparator_first_inp1_6, B0=>nx19140, B1=>nx19854);
   max_calc_reg_ans2_6 : dff port map ( Q=>max_calc_ans2_6, QB=>OPEN, D=>
      nx31021, CLK=>clk);
   max_calc_reg_ans7_6 : dff port map ( Q=>max_calc_ans7_6, QB=>OPEN, D=>
      nx31081, CLK=>clk);
   max_calc_reg_ans8_6 : dff port map ( Q=>max_calc_ans8_6, QB=>OPEN, D=>
      nx31071, CLK=>clk);
   max_calc_reg_comparator_first_inp1_6 : dff port map ( Q=>
      max_calc_comparator_first_inp1_6, QB=>OPEN, D=>nx31061, CLK=>clk);
   max_calc_reg_ans1_6 : dff port map ( Q=>max_calc_ans1_6, QB=>OPEN, D=>
      nx31031, CLK=>clk);
   max_calc_reg_ans6_6 : dff port map ( Q=>max_calc_ans6_6, QB=>OPEN, D=>
      nx31041, CLK=>clk);
   max_calc_reg_ans5_6 : dff port map ( Q=>max_calc_ans5_6, QB=>OPEN, D=>
      nx31051, CLK=>clk);
   max_calc_reg_comparator_first_inp2_6 : dff port map ( Q=>
      max_calc_comparator_first_inp2_6, QB=>nx40588, D=>nx31091, CLK=>clk);
   ix19855 : oai22 port map ( Y=>nx19854, A0=>nx40624, A1=>nx40659, B0=>
      max_calc_comparator_first_inp2_5, B1=>nx40656);
   max_calc_reg_comparator_first_inp2_5 : dff port map ( Q=>
      max_calc_comparator_first_inp2_5, QB=>OPEN, D=>nx31171, CLK=>clk);
   max_calc_reg_ans2_5 : dff port map ( Q=>max_calc_ans2_5, QB=>OPEN, D=>
      nx31101, CLK=>clk);
   max_calc_reg_ans7_5 : dff port map ( Q=>max_calc_ans7_5, QB=>OPEN, D=>
      nx31161, CLK=>clk);
   max_calc_reg_ans8_5 : dff port map ( Q=>max_calc_ans8_5, QB=>OPEN, D=>
      nx31151, CLK=>clk);
   max_calc_reg_comparator_first_inp1_5 : dff port map ( Q=>
      max_calc_comparator_first_inp1_5, QB=>nx40656, D=>nx31141, CLK=>clk);
   max_calc_reg_ans1_5 : dff port map ( Q=>max_calc_ans1_5, QB=>OPEN, D=>
      nx31111, CLK=>clk);
   max_calc_reg_ans6_5 : dff port map ( Q=>max_calc_ans6_5, QB=>OPEN, D=>
      nx31121, CLK=>clk);
   max_calc_reg_ans5_5 : dff port map ( Q=>max_calc_ans5_5, QB=>OPEN, D=>
      nx31131, CLK=>clk);
   ix40660 : aoi22 port map ( Y=>nx40659, A0=>nx40661, A1=>
      max_calc_comparator_first_inp1_4, B0=>nx19384, B1=>nx19838);
   max_calc_reg_ans2_4 : dff port map ( Q=>max_calc_ans2_4, QB=>OPEN, D=>
      nx31181, CLK=>clk);
   max_calc_reg_ans7_4 : dff port map ( Q=>max_calc_ans7_4, QB=>OPEN, D=>
      nx31241, CLK=>clk);
   max_calc_reg_ans8_4 : dff port map ( Q=>max_calc_ans8_4, QB=>OPEN, D=>
      nx31231, CLK=>clk);
   max_calc_reg_comparator_first_inp1_4 : dff port map ( Q=>
      max_calc_comparator_first_inp1_4, QB=>OPEN, D=>nx31221, CLK=>clk);
   max_calc_reg_ans1_4 : dff port map ( Q=>max_calc_ans1_4, QB=>OPEN, D=>
      nx31191, CLK=>clk);
   max_calc_reg_ans6_4 : dff port map ( Q=>max_calc_ans6_4, QB=>OPEN, D=>
      nx31201, CLK=>clk);
   max_calc_reg_ans5_4 : dff port map ( Q=>max_calc_ans5_4, QB=>OPEN, D=>
      nx31211, CLK=>clk);
   max_calc_reg_comparator_first_inp2_4 : dff port map ( Q=>
      max_calc_comparator_first_inp2_4, QB=>nx40661, D=>nx31251, CLK=>clk);
   ix19839 : oai22 port map ( Y=>nx19838, A0=>nx40697, A1=>nx40732, B0=>
      max_calc_comparator_first_inp2_3, B1=>nx40729);
   max_calc_reg_comparator_first_inp2_3 : dff port map ( Q=>
      max_calc_comparator_first_inp2_3, QB=>OPEN, D=>nx31331, CLK=>clk);
   max_calc_reg_ans2_3 : dff port map ( Q=>max_calc_ans2_3, QB=>OPEN, D=>
      nx31261, CLK=>clk);
   max_calc_reg_ans7_3 : dff port map ( Q=>max_calc_ans7_3, QB=>OPEN, D=>
      nx31321, CLK=>clk);
   max_calc_reg_ans8_3 : dff port map ( Q=>max_calc_ans8_3, QB=>OPEN, D=>
      nx31311, CLK=>clk);
   max_calc_reg_comparator_first_inp1_3 : dff port map ( Q=>
      max_calc_comparator_first_inp1_3, QB=>nx40729, D=>nx31301, CLK=>clk);
   max_calc_reg_ans1_3 : dff port map ( Q=>max_calc_ans1_3, QB=>OPEN, D=>
      nx31271, CLK=>clk);
   max_calc_reg_ans6_3 : dff port map ( Q=>max_calc_ans6_3, QB=>OPEN, D=>
      nx31281, CLK=>clk);
   max_calc_reg_ans5_3 : dff port map ( Q=>max_calc_ans5_3, QB=>OPEN, D=>
      nx31291, CLK=>clk);
   ix40733 : aoi22 port map ( Y=>nx40732, A0=>nx40734, A1=>
      max_calc_comparator_first_inp1_2, B0=>nx19628, B1=>nx19822);
   max_calc_reg_ans2_2 : dff port map ( Q=>max_calc_ans2_2, QB=>OPEN, D=>
      nx31341, CLK=>clk);
   max_calc_reg_ans7_2 : dff port map ( Q=>max_calc_ans7_2, QB=>OPEN, D=>
      nx31401, CLK=>clk);
   max_calc_reg_ans8_2 : dff port map ( Q=>max_calc_ans8_2, QB=>OPEN, D=>
      nx31391, CLK=>clk);
   max_calc_reg_comparator_first_inp1_2 : dff port map ( Q=>
      max_calc_comparator_first_inp1_2, QB=>OPEN, D=>nx31381, CLK=>clk);
   max_calc_reg_ans1_2 : dff port map ( Q=>max_calc_ans1_2, QB=>OPEN, D=>
      nx31351, CLK=>clk);
   max_calc_reg_ans6_2 : dff port map ( Q=>max_calc_ans6_2, QB=>OPEN, D=>
      nx31361, CLK=>clk);
   max_calc_reg_ans5_2 : dff port map ( Q=>max_calc_ans5_2, QB=>OPEN, D=>
      nx31371, CLK=>clk);
   max_calc_reg_comparator_first_inp2_2 : dff port map ( Q=>
      max_calc_comparator_first_inp2_2, QB=>nx40734, D=>nx31411, CLK=>clk);
   ix19823 : oai21 port map ( Y=>nx19822, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx40800, B0=>nx40803);
   max_calc_reg_comparator_first_inp2_1 : dff port map ( Q=>
      max_calc_comparator_first_inp2_1, QB=>OPEN, D=>nx31491, CLK=>clk);
   max_calc_reg_ans2_1 : dff port map ( Q=>max_calc_ans2_1, QB=>OPEN, D=>
      nx31421, CLK=>clk);
   max_calc_reg_ans7_1 : dff port map ( Q=>max_calc_ans7_1, QB=>OPEN, D=>
      nx31481, CLK=>clk);
   max_calc_reg_ans8_1 : dff port map ( Q=>max_calc_ans8_1, QB=>OPEN, D=>
      nx31471, CLK=>clk);
   max_calc_reg_comparator_first_inp1_1 : dff port map ( Q=>
      max_calc_comparator_first_inp1_1, QB=>nx40800, D=>nx31461, CLK=>clk);
   max_calc_reg_ans1_1 : dff port map ( Q=>max_calc_ans1_1, QB=>OPEN, D=>
      nx31431, CLK=>clk);
   max_calc_reg_ans6_1 : dff port map ( Q=>max_calc_ans6_1, QB=>OPEN, D=>
      nx31441, CLK=>clk);
   max_calc_reg_ans5_1 : dff port map ( Q=>max_calc_ans5_1, QB=>OPEN, D=>
      nx31451, CLK=>clk);
   ix40804 : oai21 port map ( Y=>nx40803, A0=>nx40805, A1=>
      max_calc_comparator_first_inp1_0, B0=>nx19750);
   max_calc_reg_ans2_0 : dff port map ( Q=>max_calc_ans2_0, QB=>OPEN, D=>
      nx31501, CLK=>clk);
   max_calc_reg_ans7_0 : dff port map ( Q=>max_calc_ans7_0, QB=>OPEN, D=>
      nx31521, CLK=>clk);
   max_calc_reg_ans8_0 : dff port map ( Q=>max_calc_ans8_0, QB=>OPEN, D=>
      nx31511, CLK=>clk);
   max_calc_reg_comparator_first_inp1_0 : dff port map ( Q=>
      max_calc_comparator_first_inp1_0, QB=>OPEN, D=>nx22881, CLK=>clk);
   max_calc_reg_ans1_0 : dff port map ( Q=>max_calc_ans1_0, QB=>OPEN, D=>
      nx20831, CLK=>clk);
   max_calc_reg_ans6_0 : dff port map ( Q=>max_calc_ans6_0, QB=>OPEN, D=>
      nx20841, CLK=>clk);
   max_calc_reg_ans5_0 : dff port map ( Q=>max_calc_ans5_0, QB=>OPEN, D=>
      nx22871, CLK=>clk);
   max_calc_reg_comparator_first_inp2_0 : dff port map ( Q=>
      max_calc_comparator_first_inp2_0, QB=>nx40805, D=>nx31531, CLK=>clk);
   ix20113 : xnor2 port map ( Y=>nx20112, A0=>
      max_calc_comparator_first_inp2_15, A1=>
      max_calc_comparator_first_inp1_15);
   max_calc_reg_comparator_first_inp2_15 : dff port map ( Q=>
      max_calc_comparator_first_inp2_15, QB=>OPEN, D=>nx31651, CLK=>clk);
   lat_label_2_input_15 : latch port map ( Q=>label_2_input_15, D=>nx19948, 
      CLK=>nx41705);
   reg_label_2_input_state_machine_15 : dffr port map ( Q=>
      label_2_input_state_machine_15, QB=>OPEN, D=>nx31541, CLK=>clk, R=>rst
   );
   ix19945 : xnor2 port map ( Y=>nx19944, A0=>nx40853, A1=>nx19942);
   ix40854 : aoi22 port map ( Y=>nx40853, A0=>label_2_output_14, A1=>
      booth_booth_integration_output_1_26, B0=>nx7294, B1=>nx7296);
   labelsregfile_label2_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_2_output_15, QB=>nx40857, D=>nx31551, CLK=>clk, R=>rst);
   max_calc_reg_ans2_15 : dff port map ( Q=>max_calc_ans2_15, QB=>OPEN, D=>
      nx31561, CLK=>clk);
   max_calc_reg_ans7_15 : dff port map ( Q=>max_calc_ans7_15, QB=>OPEN, D=>
      nx31641, CLK=>clk);
   max_calc_reg_ans8_15 : dff port map ( Q=>max_calc_ans8_15, QB=>OPEN, D=>
      nx31631, CLK=>clk);
   max_calc_reg_answer_13 : dffr port map ( Q=>max_calc_answer_13, QB=>OPEN, 
      D=>nx31791, CLK=>clk, R=>rst);
   ix40880 : xnor2 port map ( Y=>nx40879, A0=>nx42205, A1=>
      label_10_output_12);
   max_calc_reg_answer_12 : dffr port map ( Q=>max_calc_answer_12, QB=>OPEN, 
      D=>nx31781, CLK=>clk, R=>rst);
   ix20817 : nand04 port map ( Y=>nx20816, A0=>nx40885, A1=>nx40890, A2=>
      nx40895, A3=>nx40900);
   max_calc_reg_answer_11 : dffr port map ( Q=>max_calc_answer_11, QB=>OPEN, 
      D=>nx31771, CLK=>clk, R=>rst);
   ix40891 : xnor2 port map ( Y=>nx40890, A0=>nx42197, A1=>
      label_10_output_10);
   max_calc_reg_answer_10 : dffr port map ( Q=>max_calc_answer_10, QB=>OPEN, 
      D=>nx31761, CLK=>clk, R=>rst);
   max_calc_reg_answer_9 : dffr port map ( Q=>max_calc_answer_9, QB=>OPEN, D
      =>nx31751, CLK=>clk, R=>rst);
   ix40901 : xnor2 port map ( Y=>nx40900, A0=>nx42189, A1=>label_10_output_8
   );
   max_calc_reg_answer_8 : dffr port map ( Q=>max_calc_answer_8, QB=>OPEN, D
      =>nx31741, CLK=>clk, R=>rst);
   ix20801 : nand04 port map ( Y=>nx20800, A0=>nx40906, A1=>nx40911, A2=>
      nx40916, A3=>nx40921);
   max_calc_reg_answer_7 : dffr port map ( Q=>max_calc_answer_7, QB=>OPEN, D
      =>nx31731, CLK=>clk, R=>rst);
   ix40912 : xnor2 port map ( Y=>nx40911, A0=>nx42181, A1=>label_10_output_6
   );
   max_calc_reg_answer_6 : dffr port map ( Q=>max_calc_answer_6, QB=>OPEN, D
      =>nx31721, CLK=>clk, R=>rst);
   max_calc_reg_answer_5 : dffr port map ( Q=>max_calc_answer_5, QB=>OPEN, D
      =>nx31711, CLK=>clk, R=>rst);
   ix40922 : xnor2 port map ( Y=>nx40921, A0=>nx42173, A1=>label_10_output_4
   );
   max_calc_reg_answer_4 : dffr port map ( Q=>max_calc_answer_4, QB=>OPEN, D
      =>nx31701, CLK=>clk, R=>rst);
   ix20787 : nand04 port map ( Y=>nx20786, A0=>nx40927, A1=>nx40932, A2=>
      nx40937, A3=>nx40942);
   max_calc_reg_answer_3 : dffr port map ( Q=>max_calc_answer_3, QB=>OPEN, D
      =>nx31691, CLK=>clk, R=>rst);
   ix40933 : xnor2 port map ( Y=>nx40932, A0=>nx42165, A1=>label_10_output_2
   );
   max_calc_reg_answer_2 : dffr port map ( Q=>max_calc_answer_2, QB=>OPEN, D
      =>nx31681, CLK=>clk, R=>rst);
   max_calc_reg_answer_1 : dffr port map ( Q=>max_calc_answer_1, QB=>OPEN, D
      =>nx31671, CLK=>clk, R=>rst);
   ix40943 : xnor2 port map ( Y=>nx40942, A0=>nx41531, A1=>label_10_output_0
   );
   max_calc_reg_answer_0 : dffr port map ( Q=>max_calc_answer_0, QB=>OPEN, D
      =>nx31661, CLK=>clk, R=>rst);
   ix40948 : nor04 port map ( Y=>nx40947, A0=>nx20892, A1=>nx20878, A2=>
      nx20862, A3=>nx20848);
   ix20893 : nand04 port map ( Y=>nx20892, A0=>nx40950, A1=>nx40952, A2=>
      nx40954, A3=>nx40956);
   ix40953 : xnor2 port map ( Y=>nx40952, A0=>nx42213, A1=>label_9_output_14
   );
   ix40957 : xnor2 port map ( Y=>nx40956, A0=>nx42205, A1=>label_9_output_12
   );
   ix20879 : nand04 port map ( Y=>nx20878, A0=>nx40959, A1=>nx40961, A2=>
      nx40963, A3=>nx40965);
   ix40962 : xnor2 port map ( Y=>nx40961, A0=>nx42197, A1=>label_9_output_10
   );
   ix40966 : xnor2 port map ( Y=>nx40965, A0=>nx42189, A1=>label_9_output_8
   );
   ix20863 : nand04 port map ( Y=>nx20862, A0=>nx40968, A1=>nx40970, A2=>
      nx40972, A3=>nx40974);
   ix40971 : xnor2 port map ( Y=>nx40970, A0=>nx42181, A1=>label_9_output_6
   );
   ix40975 : xnor2 port map ( Y=>nx40974, A0=>nx42173, A1=>label_9_output_4
   );
   ix20849 : nand04 port map ( Y=>nx20848, A0=>nx40977, A1=>nx40979, A2=>
      nx40981, A3=>nx40983);
   ix40980 : xnor2 port map ( Y=>nx40979, A0=>nx42165, A1=>label_9_output_2
   );
   ix40984 : xnor2 port map ( Y=>nx40983, A0=>nx41531, A1=>label_9_output_0
   );
   max_calc_reg_ans6_15 : dff port map ( Q=>max_calc_ans6_15, QB=>OPEN, D=>
      nx31601, CLK=>clk);
   max_calc_reg_ans5_15 : dff port map ( Q=>max_calc_ans5_15, QB=>OPEN, D=>
      nx31611, CLK=>clk);
   ix40999 : xnor2 port map ( Y=>nx40998, A0=>nx42213, A1=>label_7_output_14
   );
   ix41003 : xnor2 port map ( Y=>nx41002, A0=>nx42205, A1=>label_7_output_12
   );
   ix20293 : nand04 port map ( Y=>nx20292, A0=>nx41005, A1=>nx41007, A2=>
      nx41009, A3=>nx41011);
   ix41008 : xnor2 port map ( Y=>nx41007, A0=>nx42197, A1=>label_7_output_10
   );
   ix41012 : xnor2 port map ( Y=>nx41011, A0=>nx42189, A1=>label_7_output_8
   );
   ix20277 : nand04 port map ( Y=>nx20276, A0=>nx41014, A1=>nx41016, A2=>
      nx41018, A3=>nx41020);
   ix41017 : xnor2 port map ( Y=>nx41016, A0=>nx42181, A1=>label_7_output_6
   );
   ix41021 : xnor2 port map ( Y=>nx41020, A0=>nx42173, A1=>label_7_output_4
   );
   ix20263 : nand04 port map ( Y=>nx20262, A0=>nx41023, A1=>nx41025, A2=>
      nx41027, A3=>nx41029);
   ix41026 : xnor2 port map ( Y=>nx41025, A0=>nx42165, A1=>label_7_output_2
   );
   ix41030 : xnor2 port map ( Y=>nx41029, A0=>nx41531, A1=>label_7_output_0
   );
   ix41032 : nor03_2x port map ( Y=>nx41031, A0=>nx20758, A1=>nx20664, A2=>
      nx41233);
   ix20759 : nor04 port map ( Y=>nx20758, A0=>nx41034, A1=>nx41044, A2=>
      nx41054, A3=>nx41064);
   ix41035 : nand04 port map ( Y=>nx41034, A0=>nx41036, A1=>nx41038, A2=>
      nx41040, A3=>nx41042);
   ix41037 : xnor2 port map ( Y=>nx41036, A0=>nx41531, A1=>label_6_output_0
   );
   ix41041 : xnor2 port map ( Y=>nx41040, A0=>nx42165, A1=>label_6_output_2
   );
   ix41045 : nand04 port map ( Y=>nx41044, A0=>nx41046, A1=>nx41048, A2=>
      nx41050, A3=>nx41052);
   ix41047 : xnor2 port map ( Y=>nx41046, A0=>nx42173, A1=>label_6_output_4
   );
   ix41051 : xnor2 port map ( Y=>nx41050, A0=>nx42181, A1=>label_6_output_6
   );
   ix41055 : nand04 port map ( Y=>nx41054, A0=>nx41056, A1=>nx41058, A2=>
      nx41060, A3=>nx41062);
   ix41057 : xnor2 port map ( Y=>nx41056, A0=>nx42189, A1=>label_6_output_8
   );
   ix41061 : xnor2 port map ( Y=>nx41060, A0=>nx42197, A1=>label_6_output_10
   );
   ix41065 : nand04 port map ( Y=>nx41064, A0=>nx41066, A1=>nx41068, A2=>
      nx41070, A3=>nx41072);
   ix41067 : xnor2 port map ( Y=>nx41066, A0=>nx42205, A1=>label_6_output_12
   );
   ix41071 : xnor2 port map ( Y=>nx41070, A0=>nx42213, A1=>label_6_output_14
   );
   ix41076 : nor02ii port map ( Y=>nx41075, A0=>nx41077, A1=>nx41115);
   ix41078 : nor04 port map ( Y=>nx41077, A0=>nx20492, A1=>nx20478, A2=>
      nx20462, A3=>nx20448);
   ix20493 : nand04 port map ( Y=>nx20492, A0=>nx41080, A1=>nx41082, A2=>
      nx41084, A3=>nx41086);
   ix41083 : xnor2 port map ( Y=>nx41082, A0=>nx42213, A1=>label_3_output_14
   );
   ix41087 : xnor2 port map ( Y=>nx41086, A0=>nx42205, A1=>label_3_output_12
   );
   ix20479 : nand04 port map ( Y=>nx20478, A0=>nx41089, A1=>nx41091, A2=>
      nx41093, A3=>nx41095);
   ix41092 : xnor2 port map ( Y=>nx41091, A0=>nx42197, A1=>label_3_output_10
   );
   ix41096 : xnor2 port map ( Y=>nx41095, A0=>nx42189, A1=>label_3_output_8
   );
   ix20463 : nand04 port map ( Y=>nx20462, A0=>nx41098, A1=>nx41100, A2=>
      nx41102, A3=>nx41104);
   ix41101 : xnor2 port map ( Y=>nx41100, A0=>nx42181, A1=>label_3_output_6
   );
   ix41105 : xnor2 port map ( Y=>nx41104, A0=>nx42173, A1=>label_3_output_4
   );
   ix20449 : nand04 port map ( Y=>nx20448, A0=>nx41107, A1=>nx41109, A2=>
      nx41111, A3=>nx41113);
   ix41110 : xnor2 port map ( Y=>nx41109, A0=>nx42165, A1=>label_3_output_2
   );
   ix41114 : xnor2 port map ( Y=>nx41113, A0=>nx41531, A1=>label_3_output_0
   );
   ix41116 : nor02_2x port map ( Y=>nx41115, A0=>nx20652, A1=>nx41158);
   ix20653 : nor04 port map ( Y=>nx20652, A0=>nx41118, A1=>nx41128, A2=>
      nx41138, A3=>nx41148);
   ix41119 : nand04 port map ( Y=>nx41118, A0=>nx41120, A1=>nx41122, A2=>
      nx41124, A3=>nx41126);
   ix41121 : xnor2 port map ( Y=>nx41120, A0=>nx41531, A1=>label_2_output_0
   );
   ix41125 : xnor2 port map ( Y=>nx41124, A0=>nx42165, A1=>label_2_output_2
   );
   ix41129 : nand04 port map ( Y=>nx41128, A0=>nx41130, A1=>nx41132, A2=>
      nx41134, A3=>nx41136);
   ix41131 : xnor2 port map ( Y=>nx41130, A0=>nx42173, A1=>label_2_output_4
   );
   ix41135 : xnor2 port map ( Y=>nx41134, A0=>nx42181, A1=>label_2_output_6
   );
   ix41139 : nand04 port map ( Y=>nx41138, A0=>nx41140, A1=>nx41142, A2=>
      nx41144, A3=>nx41146);
   ix41141 : xnor2 port map ( Y=>nx41140, A0=>nx42189, A1=>label_2_output_8
   );
   ix41145 : xnor2 port map ( Y=>nx41144, A0=>nx42197, A1=>label_2_output_10
   );
   ix41149 : nand04 port map ( Y=>nx41148, A0=>nx41150, A1=>nx41152, A2=>
      nx41154, A3=>nx41156);
   ix41151 : xnor2 port map ( Y=>nx41150, A0=>nx42205, A1=>label_2_output_12
   );
   ix41155 : xnor2 port map ( Y=>nx41154, A0=>nx42213, A1=>label_2_output_14
   );
   ix41159 : nor04 port map ( Y=>nx41158, A0=>nx20554, A1=>nx20540, A2=>
      nx20524, A3=>nx20510);
   ix20555 : nand04 port map ( Y=>nx20554, A0=>nx41161, A1=>nx41163, A2=>
      nx41165, A3=>nx41167);
   ix41164 : xnor2 port map ( Y=>nx41163, A0=>nx42215, A1=>label_1_output_14
   );
   ix41168 : xnor2 port map ( Y=>nx41167, A0=>nx42207, A1=>label_1_output_12
   );
   ix20541 : nand04 port map ( Y=>nx20540, A0=>nx41170, A1=>nx41172, A2=>
      nx41174, A3=>nx41176);
   ix41173 : xnor2 port map ( Y=>nx41172, A0=>nx42199, A1=>label_1_output_10
   );
   ix41177 : xnor2 port map ( Y=>nx41176, A0=>nx42191, A1=>label_1_output_8
   );
   ix20525 : nand04 port map ( Y=>nx20524, A0=>nx41179, A1=>nx41181, A2=>
      nx41183, A3=>nx41185);
   ix41182 : xnor2 port map ( Y=>nx41181, A0=>nx42183, A1=>label_1_output_6
   );
   ix41186 : xnor2 port map ( Y=>nx41185, A0=>nx42175, A1=>label_1_output_4
   );
   ix20511 : nand04 port map ( Y=>nx20510, A0=>nx41188, A1=>nx41190, A2=>
      nx41192, A3=>nx41194);
   ix41191 : xnor2 port map ( Y=>nx41190, A0=>nx42167, A1=>label_1_output_2
   );
   ix41195 : xnor2 port map ( Y=>nx41194, A0=>nx41533, A1=>label_1_output_0
   );
   ix20431 : nand04 port map ( Y=>nx20430, A0=>nx41198, A1=>nx41200, A2=>
      nx41202, A3=>nx41204);
   ix41201 : xnor2 port map ( Y=>nx41200, A0=>nx42215, A1=>label_4_output_14
   );
   ix41205 : xnor2 port map ( Y=>nx41204, A0=>nx42207, A1=>label_4_output_12
   );
   ix20417 : nand04 port map ( Y=>nx20416, A0=>nx41207, A1=>nx41209, A2=>
      nx41211, A3=>nx41213);
   ix41210 : xnor2 port map ( Y=>nx41209, A0=>nx42199, A1=>label_4_output_10
   );
   ix41214 : xnor2 port map ( Y=>nx41213, A0=>nx42191, A1=>label_4_output_8
   );
   ix20401 : nand04 port map ( Y=>nx20400, A0=>nx41216, A1=>nx41218, A2=>
      nx41220, A3=>nx41222);
   ix41219 : xnor2 port map ( Y=>nx41218, A0=>nx42183, A1=>label_4_output_6
   );
   ix41223 : xnor2 port map ( Y=>nx41222, A0=>nx42175, A1=>label_4_output_4
   );
   ix20387 : nand04 port map ( Y=>nx20386, A0=>nx41225, A1=>nx41227, A2=>
      nx41229, A3=>nx41231);
   ix41228 : xnor2 port map ( Y=>nx41227, A0=>nx42167, A1=>label_4_output_2
   );
   ix41232 : xnor2 port map ( Y=>nx41231, A0=>nx41533, A1=>label_4_output_0
   );
   ix41234 : nor04 port map ( Y=>nx41233, A0=>nx20368, A1=>nx20354, A2=>
      nx20338, A3=>nx20324);
   ix20369 : nand04 port map ( Y=>nx20368, A0=>nx41236, A1=>nx41238, A2=>
      nx41240, A3=>nx41242);
   ix41239 : xnor2 port map ( Y=>nx41238, A0=>nx42215, A1=>label_5_output_14
   );
   ix41243 : xnor2 port map ( Y=>nx41242, A0=>nx42207, A1=>label_5_output_12
   );
   ix20355 : nand04 port map ( Y=>nx20354, A0=>nx41245, A1=>nx41247, A2=>
      nx41249, A3=>nx41251);
   ix41248 : xnor2 port map ( Y=>nx41247, A0=>nx42199, A1=>label_5_output_10
   );
   ix41252 : xnor2 port map ( Y=>nx41251, A0=>nx42191, A1=>label_5_output_8
   );
   ix20339 : nand04 port map ( Y=>nx20338, A0=>nx41254, A1=>nx41256, A2=>
      nx41258, A3=>nx41260);
   ix41257 : xnor2 port map ( Y=>nx41256, A0=>nx42183, A1=>label_5_output_6
   );
   ix41261 : xnor2 port map ( Y=>nx41260, A0=>nx42175, A1=>label_5_output_4
   );
   ix20325 : nand04 port map ( Y=>nx20324, A0=>nx41263, A1=>nx41265, A2=>
      nx41267, A3=>nx41269);
   ix41266 : xnor2 port map ( Y=>nx41265, A0=>nx42167, A1=>label_5_output_2
   );
   ix41270 : xnor2 port map ( Y=>nx41269, A0=>nx41533, A1=>label_5_output_0
   );
   ix20245 : nand04 port map ( Y=>nx20244, A0=>nx41273, A1=>nx41275, A2=>
      nx41277, A3=>nx41279);
   ix41276 : xnor2 port map ( Y=>nx41275, A0=>nx42215, A1=>label_8_output_14
   );
   ix41280 : xnor2 port map ( Y=>nx41279, A0=>nx42207, A1=>label_8_output_12
   );
   ix20215 : nand04 port map ( Y=>nx20214, A0=>nx41282, A1=>nx41284, A2=>
      nx41286, A3=>nx41288);
   ix41285 : xnor2 port map ( Y=>nx41284, A0=>nx42199, A1=>label_8_output_10
   );
   ix41289 : xnor2 port map ( Y=>nx41288, A0=>nx42191, A1=>label_8_output_8
   );
   ix20183 : nand04 port map ( Y=>nx20182, A0=>nx41291, A1=>nx41293, A2=>
      nx41295, A3=>nx41297);
   ix41294 : xnor2 port map ( Y=>nx41293, A0=>nx42183, A1=>label_8_output_6
   );
   ix41298 : xnor2 port map ( Y=>nx41297, A0=>nx42175, A1=>label_8_output_4
   );
   ix20153 : nand04 port map ( Y=>nx20152, A0=>nx41300, A1=>nx41302, A2=>
      nx41304, A3=>nx41306);
   ix41303 : xnor2 port map ( Y=>nx41302, A0=>nx42167, A1=>label_8_output_2
   );
   ix41307 : xnor2 port map ( Y=>nx41306, A0=>nx41533, A1=>label_8_output_0
   );
   ix41311 : aoi32 port map ( Y=>nx41310, A0=>nx42245, A1=>nx41371, A2=>
      nx34114, B0=>nx33436, B1=>nx1758);
   ix1759 : aoi21 port map ( Y=>nx1758, A0=>nx34114, A1=>nx42245, B0=>
      nx41373);
   max_calc_reg_result_0 : dffr port map ( Q=>answer_0_EXMPLR, QB=>OPEN, D=>
      nx31841, CLK=>clk, R=>rst);
   ix31842 : mux21_ni port map ( Y=>nx31841, A0=>answer_0_EXMPLR, A1=>
      nx20988, S0=>nx20950);
   ix20989 : nand03 port map ( Y=>nx20988, A0=>nx41319, A1=>nx20558, A2=>
      nx41328);
   ix41320 : nand02 port map ( Y=>nx41319, A0=>nx40947, A1=>nx41321);
   ix41326 : nor04 port map ( Y=>nx41325, A0=>nx20244, A1=>nx20214, A2=>
      nx20182, A3=>nx20152);
   ix41329 : aoi222 port map ( Y=>nx41328, A0=>nx41077, A1=>nx41115, B0=>
      nx41233, B1=>nx41330, C0=>nx32711, C1=>nx41031);
   ix41331 : nor02ii port map ( Y=>nx41330, A0=>nx41332, A1=>nx41075);
   ix41333 : nor04 port map ( Y=>nx41332, A0=>nx20430, A1=>nx20416, A2=>
      nx20400, A3=>nx20386);
   max_calc_reg_result_1 : dffr port map ( Q=>answer_1_EXMPLR, QB=>OPEN, D=>
      nx31851, CLK=>clk, R=>rst);
   ix31852 : mux21_ni port map ( Y=>nx31851, A0=>answer_1_EXMPLR, A1=>
      nx21008, S0=>nx20950);
   ix21009 : and04 port map ( Y=>nx21008, A0=>nx20558, A1=>nx41319, A2=>
      nx21002, A3=>nx21004);
   ix21003 : oai21 port map ( Y=>nx21002, A0=>nx41332, A1=>nx41233, B0=>
      nx41075);
   ix21005 : nand02 port map ( Y=>nx21004, A0=>nx32709, A1=>nx41325);
   max_calc_reg_result_2 : dffr port map ( Q=>answer_2_EXMPLR, QB=>OPEN, D=>
      nx31861, CLK=>clk, R=>rst);
   ix31862 : mux21_ni port map ( Y=>nx31861, A0=>answer_2_EXMPLR, A1=>
      nx21016, S0=>nx20950);
   ix21017 : nor02ii port map ( Y=>nx21016, A0=>nx32709, A1=>nx41075);
   max_calc_reg_result_3 : dffr port map ( Q=>answer_3_EXMPLR, QB=>OPEN, D=>
      nx31871, CLK=>clk, R=>rst);
   ix31872 : mux21_ni port map ( Y=>nx31871, A0=>answer_3_EXMPLR, A1=>
      nx21034, S0=>nx20950);
   ix21035 : nand02 port map ( Y=>nx21034, A0=>nx41348, A1=>nx41319);
   ix41349 : mux21 port map ( Y=>nx41348, A0=>nx32709, A1=>nx33450, S0=>
      nx41321);
   reg_enable_read : dffr port map ( Q=>enable_read_EXMPLR, QB=>OPEN, D=>
      nx31881, CLK=>clk, R=>rst);
   ix31882 : mux21_ni port map ( Y=>nx31881, A0=>enable_read_EXMPLR, A1=>
      nx1612, S0=>nx21076);
   ix41355 : aoi21 port map ( Y=>nx41354, A0=>nx42887, A1=>nx41379, B0=>
      nx42865);
   ix21077 : aoi21 port map ( Y=>nx21076, A0=>nx41357, A1=>nx41362, B0=>
      nx104);
   ix41358 : oai21 port map ( Y=>nx41357, A0=>nx21062, A1=>nx42257, B0=>
      nx41360);
   ix41363 : nand03 port map ( Y=>nx41362, A0=>nx21046, A1=>nx43041, A2=>
      nx31914);
   ix20773 : inv01 port map ( Y=>nx20772, A=>nx41321);
   ix20665 : inv01 port map ( Y=>nx20664, A=>nx41330);
   ix20559 : inv01 port map ( Y=>nx20558, A=>nx41158);
   ix18053 : inv01 port map ( Y=>nx18052, A=>nx33416);
   ix18013 : inv01 port map ( Y=>nx18599, A=>nx33401);
   ix17949 : inv01 port map ( Y=>nx18597, A=>nx33386);
   ix17885 : inv01 port map ( Y=>nx18595, A=>nx33371);
   ix17821 : inv01 port map ( Y=>nx18593, A=>nx33356);
   ix17757 : inv01 port map ( Y=>nx18589, A=>nx33341);
   ix17693 : inv01 port map ( Y=>nx18585, A=>nx33326);
   ix15735 : inv01 port map ( Y=>nx15734, A=>nx39686);
   ix15695 : inv01 port map ( Y=>nx18580, A=>nx39671);
   ix15631 : inv01 port map ( Y=>nx18578, A=>nx39656);
   ix15567 : inv01 port map ( Y=>nx18576, A=>nx39641);
   ix15503 : inv01 port map ( Y=>nx18573, A=>nx39626);
   ix15439 : inv01 port map ( Y=>nx18569, A=>nx39611);
   ix15375 : inv01 port map ( Y=>nx18566, A=>nx39596);
   ix39539 : inv01 port map ( Y=>nx39538, A=>nx18563);
   ix15017 : inv01 port map ( Y=>nx15016, A=>nx39556);
   ix39544 : inv01 port map ( Y=>nx39543, A=>nx15006);
   ix39501 : inv01 port map ( Y=>nx39500, A=>nx18561);
   ix14969 : inv01 port map ( Y=>nx14968, A=>nx39559);
   ix39506 : inv01 port map ( Y=>nx39505, A=>nx14958);
   ix39465 : inv01 port map ( Y=>nx39464, A=>nx18557);
   ix14921 : inv01 port map ( Y=>nx14920, A=>nx39562);
   ix39470 : inv01 port map ( Y=>nx39469, A=>nx14910);
   ix39429 : inv01 port map ( Y=>nx39428, A=>nx18553);
   ix14873 : inv01 port map ( Y=>nx14872, A=>nx39565);
   ix39434 : inv01 port map ( Y=>nx39433, A=>nx14862);
   ix39393 : inv01 port map ( Y=>nx39392, A=>nx18549);
   ix14825 : inv01 port map ( Y=>nx14824, A=>nx39568);
   ix39398 : inv01 port map ( Y=>nx39397, A=>nx14814);
   ix39357 : inv01 port map ( Y=>nx39356, A=>nx18547);
   ix39362 : inv01 port map ( Y=>nx39361, A=>nx14766);
   ix15199 : inv01 port map ( Y=>nx18546, A=>nx39330);
   ix39327 : inv01 port map ( Y=>nx39326, A=>nx14742);
   ix39322 : inv01 port map ( Y=>nx39321, A=>nx18545);
   ix14729 : inv01 port map ( Y=>nx14728, A=>nx39571);
   ix39575 : inv01 port map ( Y=>nx39574, A=>nx14718);
   ix14419 : inv01 port map ( Y=>nx14418, A=>nx39052);
   ix14379 : inv01 port map ( Y=>nx18539, A=>nx39037);
   ix14315 : inv01 port map ( Y=>nx18535, A=>nx39022);
   ix14251 : inv01 port map ( Y=>nx18531, A=>nx39007);
   ix14187 : inv01 port map ( Y=>nx18528, A=>nx38992);
   ix14123 : inv01 port map ( Y=>nx18526, A=>nx38977);
   ix14059 : inv01 port map ( Y=>nx18524, A=>nx38962);
   ix38905 : inv01 port map ( Y=>nx38904, A=>nx18519);
   ix13701 : inv01 port map ( Y=>nx13700, A=>nx38922);
   ix38910 : inv01 port map ( Y=>nx38909, A=>nx13690);
   ix38867 : inv01 port map ( Y=>nx38866, A=>nx18515);
   ix13653 : inv01 port map ( Y=>nx13652, A=>nx38925);
   ix38872 : inv01 port map ( Y=>nx38871, A=>nx13642);
   ix38831 : inv01 port map ( Y=>nx38830, A=>nx18512);
   ix13605 : inv01 port map ( Y=>nx13604, A=>nx38928);
   ix38836 : inv01 port map ( Y=>nx38835, A=>nx13594);
   ix38795 : inv01 port map ( Y=>nx38794, A=>nx18510);
   ix13557 : inv01 port map ( Y=>nx13556, A=>nx38931);
   ix38800 : inv01 port map ( Y=>nx38799, A=>nx13546);
   ix38759 : inv01 port map ( Y=>nx38758, A=>nx18508);
   ix13509 : inv01 port map ( Y=>nx13508, A=>nx38934);
   ix38764 : inv01 port map ( Y=>nx38763, A=>nx13498);
   ix38723 : inv01 port map ( Y=>nx38722, A=>nx18505);
   ix38728 : inv01 port map ( Y=>nx38727, A=>nx13450);
   ix13883 : inv01 port map ( Y=>nx18504, A=>nx38696);
   ix38693 : inv01 port map ( Y=>nx38692, A=>nx13426);
   ix38688 : inv01 port map ( Y=>nx38687, A=>nx18503);
   ix13413 : inv01 port map ( Y=>nx13412, A=>nx38937);
   ix38941 : inv01 port map ( Y=>nx38940, A=>nx13402);
   ix13109 : inv01 port map ( Y=>nx13108, A=>nx38415);
   ix13069 : inv01 port map ( Y=>nx18499, A=>nx38400);
   ix13005 : inv01 port map ( Y=>nx18497, A=>nx38385);
   ix12941 : inv01 port map ( Y=>nx18493, A=>nx38370);
   ix12877 : inv01 port map ( Y=>nx18490, A=>nx38355);
   ix12813 : inv01 port map ( Y=>nx18488, A=>nx38340);
   ix12749 : inv01 port map ( Y=>nx18486, A=>nx38325);
   ix38268 : inv01 port map ( Y=>nx38267, A=>nx18481);
   ix12391 : inv01 port map ( Y=>nx12390, A=>nx38285);
   ix38273 : inv01 port map ( Y=>nx38272, A=>nx12380);
   ix38230 : inv01 port map ( Y=>nx38229, A=>nx18477);
   ix12343 : inv01 port map ( Y=>nx12342, A=>nx38288);
   ix38235 : inv01 port map ( Y=>nx38234, A=>nx12332);
   ix38194 : inv01 port map ( Y=>nx38193, A=>nx18475);
   ix12295 : inv01 port map ( Y=>nx12294, A=>nx38291);
   ix38199 : inv01 port map ( Y=>nx38198, A=>nx12284);
   ix38158 : inv01 port map ( Y=>nx38157, A=>nx18473);
   ix12247 : inv01 port map ( Y=>nx12246, A=>nx38294);
   ix38163 : inv01 port map ( Y=>nx38162, A=>nx12236);
   ix38122 : inv01 port map ( Y=>nx38121, A=>nx18471);
   ix12199 : inv01 port map ( Y=>nx12198, A=>nx38297);
   ix38127 : inv01 port map ( Y=>nx38126, A=>nx12188);
   ix38086 : inv01 port map ( Y=>nx38085, A=>nx18467);
   ix38091 : inv01 port map ( Y=>nx38090, A=>nx12140);
   ix12573 : inv01 port map ( Y=>nx18465, A=>nx38059);
   ix38056 : inv01 port map ( Y=>nx38055, A=>nx12116);
   ix38051 : inv01 port map ( Y=>nx38050, A=>nx18463);
   ix12103 : inv01 port map ( Y=>nx12102, A=>nx38300);
   ix38304 : inv01 port map ( Y=>nx38303, A=>nx12092);
   ix11245 : inv01 port map ( Y=>nx11244, A=>nx37536);
   ix11205 : inv01 port map ( Y=>nx18457, A=>nx37521);
   ix11141 : inv01 port map ( Y=>nx18455, A=>nx37506);
   ix11077 : inv01 port map ( Y=>nx18453, A=>nx37491);
   ix11013 : inv01 port map ( Y=>nx18449, A=>nx37476);
   ix10949 : inv01 port map ( Y=>nx18445, A=>nx37461);
   ix10885 : inv01 port map ( Y=>nx18443, A=>nx37446);
   ix37389 : inv01 port map ( Y=>nx37388, A=>nx18440);
   ix10527 : inv01 port map ( Y=>nx10526, A=>nx37406);
   ix37394 : inv01 port map ( Y=>nx37393, A=>nx10516);
   ix37351 : inv01 port map ( Y=>nx37350, A=>nx18437);
   ix10479 : inv01 port map ( Y=>nx10478, A=>nx37409);
   ix37356 : inv01 port map ( Y=>nx37355, A=>nx10468);
   ix37315 : inv01 port map ( Y=>nx37314, A=>nx18433);
   ix10431 : inv01 port map ( Y=>nx10430, A=>nx37412);
   ix37320 : inv01 port map ( Y=>nx37319, A=>nx10420);
   ix37279 : inv01 port map ( Y=>nx37278, A=>nx18429);
   ix10383 : inv01 port map ( Y=>nx10382, A=>nx37415);
   ix37284 : inv01 port map ( Y=>nx37283, A=>nx10372);
   ix37243 : inv01 port map ( Y=>nx37242, A=>nx18426);
   ix10335 : inv01 port map ( Y=>nx10334, A=>nx37418);
   ix37248 : inv01 port map ( Y=>nx37247, A=>nx10324);
   ix37207 : inv01 port map ( Y=>nx37206, A=>nx18424);
   ix37212 : inv01 port map ( Y=>nx37211, A=>nx10276);
   ix10709 : inv01 port map ( Y=>nx18423, A=>nx37180);
   ix37177 : inv01 port map ( Y=>nx37176, A=>nx10252);
   ix37172 : inv01 port map ( Y=>nx37171, A=>nx18422);
   ix10239 : inv01 port map ( Y=>nx10238, A=>nx37421);
   ix37425 : inv01 port map ( Y=>nx37424, A=>nx10228);
   ix9927 : inv01 port map ( Y=>nx9926, A=>nx36900);
   ix9887 : inv01 port map ( Y=>nx18415, A=>nx36885);
   ix9823 : inv01 port map ( Y=>nx18411, A=>nx36870);
   ix9759 : inv01 port map ( Y=>nx18407, A=>nx36855);
   ix9695 : inv01 port map ( Y=>nx18405, A=>nx36840);
   ix9631 : inv01 port map ( Y=>nx18403, A=>nx36825);
   ix9567 : inv01 port map ( Y=>nx18401, A=>nx36810);
   ix36753 : inv01 port map ( Y=>nx36752, A=>nx18395);
   ix9209 : inv01 port map ( Y=>nx9208, A=>nx36770);
   ix36758 : inv01 port map ( Y=>nx36757, A=>nx9198);
   ix36715 : inv01 port map ( Y=>nx36714, A=>nx18391);
   ix9161 : inv01 port map ( Y=>nx9160, A=>nx36773);
   ix36720 : inv01 port map ( Y=>nx36719, A=>nx9150);
   ix36679 : inv01 port map ( Y=>nx36678, A=>nx18389);
   ix9113 : inv01 port map ( Y=>nx9112, A=>nx36776);
   ix36684 : inv01 port map ( Y=>nx36683, A=>nx9102);
   ix36643 : inv01 port map ( Y=>nx36642, A=>nx18387);
   ix9065 : inv01 port map ( Y=>nx9064, A=>nx36779);
   ix36648 : inv01 port map ( Y=>nx36647, A=>nx9054);
   ix36607 : inv01 port map ( Y=>nx36606, A=>nx18385);
   ix9017 : inv01 port map ( Y=>nx9016, A=>nx36782);
   ix36612 : inv01 port map ( Y=>nx36611, A=>nx9006);
   ix36571 : inv01 port map ( Y=>nx36570, A=>nx18382);
   ix36576 : inv01 port map ( Y=>nx36575, A=>nx8958);
   ix9391 : inv01 port map ( Y=>nx18381, A=>nx36544);
   ix36541 : inv01 port map ( Y=>nx36540, A=>nx8934);
   ix36536 : inv01 port map ( Y=>nx36535, A=>nx18380);
   ix8921 : inv01 port map ( Y=>nx8920, A=>nx36785);
   ix36789 : inv01 port map ( Y=>nx36788, A=>nx8910);
   ix8607 : inv01 port map ( Y=>nx8606, A=>nx36263);
   ix8567 : inv01 port map ( Y=>nx18376, A=>nx36248);
   ix8503 : inv01 port map ( Y=>nx18373, A=>nx36233);
   ix8439 : inv01 port map ( Y=>nx18369, A=>nx36218);
   ix8375 : inv01 port map ( Y=>nx18367, A=>nx36203);
   ix8311 : inv01 port map ( Y=>nx18365, A=>nx36188);
   ix8247 : inv01 port map ( Y=>nx18363, A=>nx36173);
   ix36116 : inv01 port map ( Y=>nx36115, A=>nx18357);
   ix7889 : inv01 port map ( Y=>nx7888, A=>nx36133);
   ix36121 : inv01 port map ( Y=>nx36120, A=>nx7878);
   ix36078 : inv01 port map ( Y=>nx36077, A=>nx18354);
   ix7841 : inv01 port map ( Y=>nx7840, A=>nx36136);
   ix36083 : inv01 port map ( Y=>nx36082, A=>nx7830);
   ix36042 : inv01 port map ( Y=>nx36041, A=>nx18352);
   ix7793 : inv01 port map ( Y=>nx7792, A=>nx36139);
   ix36047 : inv01 port map ( Y=>nx36046, A=>nx7782);
   ix36006 : inv01 port map ( Y=>nx36005, A=>nx18350);
   ix7745 : inv01 port map ( Y=>nx7744, A=>nx36142);
   ix36011 : inv01 port map ( Y=>nx36010, A=>nx7734);
   ix35970 : inv01 port map ( Y=>nx35969, A=>nx18347);
   ix7697 : inv01 port map ( Y=>nx7696, A=>nx36145);
   ix35975 : inv01 port map ( Y=>nx35974, A=>nx7686);
   ix35934 : inv01 port map ( Y=>nx35933, A=>nx18343);
   ix35939 : inv01 port map ( Y=>nx35938, A=>nx7638);
   ix8071 : inv01 port map ( Y=>nx18341, A=>nx35907);
   ix35904 : inv01 port map ( Y=>nx35903, A=>nx7614);
   ix35899 : inv01 port map ( Y=>nx35898, A=>nx18339);
   ix7601 : inv01 port map ( Y=>nx7600, A=>nx36148);
   ix36152 : inv01 port map ( Y=>nx36151, A=>nx7590);
   ix7297 : inv01 port map ( Y=>nx7296, A=>nx35625);
   ix7257 : inv01 port map ( Y=>nx18334, A=>nx35610);
   ix7193 : inv01 port map ( Y=>nx18332, A=>nx35595);
   ix7129 : inv01 port map ( Y=>nx18329, A=>nx35580);
   ix7065 : inv01 port map ( Y=>nx18325, A=>nx35565);
   ix7001 : inv01 port map ( Y=>nx18322, A=>nx35550);
   ix6937 : inv01 port map ( Y=>nx18320, A=>nx35535);
   ix35478 : inv01 port map ( Y=>nx35477, A=>nx18317);
   ix6579 : inv01 port map ( Y=>nx6578, A=>nx35495);
   ix35483 : inv01 port map ( Y=>nx35482, A=>nx6568);
   ix35440 : inv01 port map ( Y=>nx35439, A=>nx18313);
   ix6531 : inv01 port map ( Y=>nx6530, A=>nx35498);
   ix35445 : inv01 port map ( Y=>nx35444, A=>nx6520);
   ix35404 : inv01 port map ( Y=>nx35403, A=>nx18309);
   ix6483 : inv01 port map ( Y=>nx6482, A=>nx35501);
   ix35409 : inv01 port map ( Y=>nx35408, A=>nx6472);
   ix35368 : inv01 port map ( Y=>nx35367, A=>nx18305);
   ix6435 : inv01 port map ( Y=>nx6434, A=>nx35504);
   ix35373 : inv01 port map ( Y=>nx35372, A=>nx6424);
   ix35332 : inv01 port map ( Y=>nx35331, A=>nx18303);
   ix6387 : inv01 port map ( Y=>nx6386, A=>nx35507);
   ix35337 : inv01 port map ( Y=>nx35336, A=>nx6376);
   ix35296 : inv01 port map ( Y=>nx35295, A=>nx18301);
   ix35301 : inv01 port map ( Y=>nx35300, A=>nx6328);
   ix6761 : inv01 port map ( Y=>nx18300, A=>nx35269);
   ix35266 : inv01 port map ( Y=>nx35265, A=>nx6304);
   ix35261 : inv01 port map ( Y=>nx35260, A=>nx18299);
   ix6291 : inv01 port map ( Y=>nx6290, A=>nx35510);
   ix35514 : inv01 port map ( Y=>nx35513, A=>nx6280);
   ix5507 : inv01 port map ( Y=>nx5506, A=>nx34755);
   ix5467 : inv01 port map ( Y=>nx18291, A=>nx34740);
   ix5403 : inv01 port map ( Y=>nx18287, A=>nx34725);
   ix5339 : inv01 port map ( Y=>nx18284, A=>nx34710);
   ix5275 : inv01 port map ( Y=>nx18282, A=>nx34695);
   ix5211 : inv01 port map ( Y=>nx18280, A=>nx34680);
   ix5147 : inv01 port map ( Y=>nx18277, A=>nx34665);
   ix5057 : inv01 port map ( Y=>nx5056, A=>nx34090);
   ix5017 : inv01 port map ( Y=>nx18271, A=>nx34075);
   ix4953 : inv01 port map ( Y=>nx18268, A=>nx34060);
   ix4889 : inv01 port map ( Y=>nx18266, A=>nx34045);
   ix4825 : inv01 port map ( Y=>nx18264, A=>nx34030);
   ix4761 : inv01 port map ( Y=>nx18261, A=>nx34015);
   ix4697 : inv01 port map ( Y=>nx18259, A=>nx34000);
   ix33943 : inv01 port map ( Y=>nx33942, A=>nx18256);
   ix4339 : inv01 port map ( Y=>nx4338, A=>nx33960);
   ix33948 : inv01 port map ( Y=>nx33947, A=>nx4328);
   ix33905 : inv01 port map ( Y=>nx33904, A=>nx18254);
   ix4291 : inv01 port map ( Y=>nx4290, A=>nx33963);
   ix33910 : inv01 port map ( Y=>nx33909, A=>nx4280);
   ix33869 : inv01 port map ( Y=>nx33868, A=>nx18251);
   ix4243 : inv01 port map ( Y=>nx4242, A=>nx33966);
   ix33874 : inv01 port map ( Y=>nx33873, A=>nx4232);
   ix33833 : inv01 port map ( Y=>nx33832, A=>nx18247);
   ix4195 : inv01 port map ( Y=>nx4194, A=>nx33969);
   ix33838 : inv01 port map ( Y=>nx33837, A=>nx4184);
   ix33797 : inv01 port map ( Y=>nx33796, A=>nx18245);
   ix4147 : inv01 port map ( Y=>nx4146, A=>nx33972);
   ix33802 : inv01 port map ( Y=>nx33801, A=>nx4136);
   ix33761 : inv01 port map ( Y=>nx33760, A=>nx18243);
   ix33766 : inv01 port map ( Y=>nx33765, A=>nx4088);
   ix4521 : inv01 port map ( Y=>nx18242, A=>nx33734);
   ix33731 : inv01 port map ( Y=>nx33730, A=>nx4064);
   ix33726 : inv01 port map ( Y=>nx33725, A=>nx18241);
   ix4051 : inv01 port map ( Y=>nx4050, A=>nx33975);
   ix33979 : inv01 port map ( Y=>nx33978, A=>nx4040);
   ix34608 : inv01 port map ( Y=>nx34607, A=>nx18235);
   ix3459 : inv01 port map ( Y=>nx3458, A=>nx34625);
   ix34613 : inv01 port map ( Y=>nx34612, A=>nx3448);
   ix34570 : inv01 port map ( Y=>nx34569, A=>nx18232);
   ix3411 : inv01 port map ( Y=>nx3410, A=>nx34628);
   ix34575 : inv01 port map ( Y=>nx34574, A=>nx3400);
   ix34534 : inv01 port map ( Y=>nx34533, A=>nx18230);
   ix3363 : inv01 port map ( Y=>nx3362, A=>nx34631);
   ix34539 : inv01 port map ( Y=>nx34538, A=>nx3352);
   ix34498 : inv01 port map ( Y=>nx34497, A=>nx18228);
   ix3315 : inv01 port map ( Y=>nx3314, A=>nx34634);
   ix34503 : inv01 port map ( Y=>nx34502, A=>nx3304);
   ix34462 : inv01 port map ( Y=>nx34461, A=>nx18225);
   ix3267 : inv01 port map ( Y=>nx3266, A=>nx34637);
   ix34467 : inv01 port map ( Y=>nx34466, A=>nx3256);
   ix34426 : inv01 port map ( Y=>nx34425, A=>nx18221);
   ix34431 : inv01 port map ( Y=>nx34430, A=>nx3208);
   ix3641 : inv01 port map ( Y=>nx18219, A=>nx34399);
   ix34396 : inv01 port map ( Y=>nx34395, A=>nx3184);
   ix34391 : inv01 port map ( Y=>nx34390, A=>nx18217);
   ix3171 : inv01 port map ( Y=>nx3170, A=>nx34640);
   ix34644 : inv01 port map ( Y=>nx34643, A=>nx3160);
   ix33243 : inv01 port map ( Y=>nx33242, A=>nx18212);
   ix2517 : inv01 port map ( Y=>nx2516, A=>nx33258);
   ix33248 : inv01 port map ( Y=>nx33247, A=>nx2506);
   ix33207 : inv01 port map ( Y=>nx33206, A=>nx18210);
   ix2469 : inv01 port map ( Y=>nx2468, A=>nx33261);
   ix33212 : inv01 port map ( Y=>nx33211, A=>nx2458);
   ix33173 : inv01 port map ( Y=>nx33172, A=>nx18207);
   ix2421 : inv01 port map ( Y=>nx2420, A=>nx33264);
   ix33178 : inv01 port map ( Y=>nx33177, A=>nx2410);
   ix33139 : inv01 port map ( Y=>nx33138, A=>nx18203);
   ix2373 : inv01 port map ( Y=>nx2372, A=>nx33267);
   ix33144 : inv01 port map ( Y=>nx33143, A=>nx2362);
   ix33105 : inv01 port map ( Y=>nx33104, A=>nx18200);
   ix2325 : inv01 port map ( Y=>nx2324, A=>nx33270);
   ix33110 : inv01 port map ( Y=>nx33109, A=>nx2314);
   ix33071 : inv01 port map ( Y=>nx33070, A=>nx18198);
   ix33076 : inv01 port map ( Y=>nx33075, A=>nx2266);
   ix2699 : inv01 port map ( Y=>nx18197, A=>nx33044);
   ix33043 : inv01 port map ( Y=>nx33042, A=>nx2242);
   ix33038 : inv01 port map ( Y=>nx33037, A=>nx18196);
   ix2229 : inv01 port map ( Y=>nx2228, A=>nx33273);
   ix33277 : inv01 port map ( Y=>nx33276, A=>nx2218);
   ix32706 : inv01 port map ( Y=>nx32705, A=>nx18191);
   ix1805 : inv01 port map ( Y=>nx18187, A=>nx34114);
   ix1715 : inv01 port map ( Y=>nx1714, A=>nx33444);
   ix1477 : inv01 port map ( Y=>nx18181, A=>nx32619);
   ix1403 : inv01 port map ( Y=>nx1402, A=>nx32585);
   ix1325 : inv01 port map ( Y=>nx18179, A=>nx32544);
   ix1251 : inv01 port map ( Y=>nx1250, A=>nx32510);
   ix1175 : inv01 port map ( Y=>nx18177, A=>nx32470);
   ix1101 : inv01 port map ( Y=>nx1100, A=>nx32436);
   ix1021 : inv01 port map ( Y=>nx18173, A=>nx32395);
   ix947 : inv01 port map ( Y=>nx946, A=>nx32361);
   ix871 : inv01 port map ( Y=>nx18169, A=>nx32321);
   ix797 : inv01 port map ( Y=>nx796, A=>nx32287);
   ix719 : inv01 port map ( Y=>nx18165, A=>nx32246);
   ix645 : inv01 port map ( Y=>nx644, A=>nx32212);
   ix565 : inv01 port map ( Y=>nx18162, A=>nx31946);
   ix509 : inv01 port map ( Y=>nx18161, A=>nx32148);
   ix361 : inv01 port map ( Y=>nx360, A=>nx32085);
   ix33300 : inv01 port map ( Y=>nx33299, A=>nx18159);
   ix105 : inv01 port map ( Y=>nx104, A=>nx31957);
   ix31971 : inv01 port map ( Y=>nx31970, A=>nx36);
   ix41361 : inv01 port map ( Y=>nx41360, A=>nx18153);
   ix32690 : inv01 port map ( Y=>nx32689, A=>nx18146);
   ix41370 : inv02 port map ( Y=>nx41371, A=>nx33429);
   ix41372 : inv02 port map ( Y=>nx41373, A=>nx42925);
   ix41374 : inv02 port map ( Y=>nx41375, A=>nx42257);
   ix41376 : inv02 port map ( Y=>nx41377, A=>nx42257);
   ix41378 : inv02 port map ( Y=>nx41379, A=>nx42257);
   ix41380 : inv02 port map ( Y=>nx41381, A=>nx31926);
   ix41382 : inv02 port map ( Y=>nx41383, A=>nx31930);
   ix41384 : inv02 port map ( Y=>nx41385, A=>nx42883);
   ix41386 : inv02 port map ( Y=>nx41387, A=>nx42283);
   ix41388 : inv02 port map ( Y=>nx41389, A=>nx42283);
   ix41390 : inv02 port map ( Y=>nx41391, A=>nx43041);
   ix41396 : inv02 port map ( Y=>nx41397, A=>nx43041);
   ix41404 : inv02 port map ( Y=>nx41405, A=>nx31972);
   ix41406 : inv02 port map ( Y=>nx41407, A=>nx42887);
   ix41408 : inv01 port map ( Y=>nx41409, A=>nx43103);
   ix41410 : inv01 port map ( Y=>nx41411, A=>nx43103);
   ix41412 : inv04 port map ( Y=>nx41413, A=>nx43097);
   ix41414 : inv04 port map ( Y=>nx41415, A=>nx43097);
   ix41416 : inv04 port map ( Y=>nx41417, A=>nx43097);
   ix41418 : inv04 port map ( Y=>nx41419, A=>nx43097);
   ix41420 : inv02 port map ( Y=>nx41421, A=>nx43055);
   ix41424 : inv02 port map ( Y=>nx41425, A=>nx43055);
   ix41428 : inv02 port map ( Y=>nx41429, A=>nx43061);
   ix41434 : inv02 port map ( Y=>nx41435, A=>nx43061);
   ix41438 : inv02 port map ( Y=>nx41439, A=>nx43061);
   ix41442 : inv02 port map ( Y=>nx41443, A=>nx43073);
   ix41446 : inv02 port map ( Y=>nx41447, A=>nx43073);
   ix41452 : inv02 port map ( Y=>nx41453, A=>nx43073);
   ix41456 : inv02 port map ( Y=>nx41457, A=>nx43085);
   ix41460 : inv02 port map ( Y=>nx41461, A=>nx43085);
   ix41468 : inv02 port map ( Y=>nx41469, A=>ready_signal);
   ix41470 : inv02 port map ( Y=>nx41471, A=>nx42789);
   ix41472 : inv02 port map ( Y=>nx41473, A=>nx42789);
   ix41474 : inv02 port map ( Y=>nx41475, A=>nx42789);
   ix41476 : inv02 port map ( Y=>nx41477, A=>nx42789);
   ix41478 : inv02 port map ( Y=>nx41479, A=>nx42789);
   ix41480 : inv02 port map ( Y=>nx41481, A=>nx42789);
   ix41482 : inv02 port map ( Y=>nx41483, A=>nx42791);
   ix41484 : inv02 port map ( Y=>nx41485, A=>nx42791);
   ix41486 : inv02 port map ( Y=>nx41487, A=>nx42791);
   ix41488 : inv02 port map ( Y=>nx41489, A=>nx42791);
   ix41490 : inv02 port map ( Y=>nx41491, A=>nx42791);
   ix41492 : inv02 port map ( Y=>nx41493, A=>nx42791);
   ix41494 : inv02 port map ( Y=>nx41495, A=>nx42791);
   ix41496 : inv02 port map ( Y=>nx41497, A=>nx42793);
   ix41498 : inv02 port map ( Y=>nx41499, A=>nx42793);
   ix41500 : inv02 port map ( Y=>nx41501, A=>nx42793);
   ix41502 : inv02 port map ( Y=>nx41503, A=>nx42793);
   ix41504 : inv02 port map ( Y=>nx41505, A=>nx42793);
   ix41514 : inv02 port map ( Y=>nx41515, A=>nx42965);
   ix41522 : inv02 port map ( Y=>nx41523, A=>nx41521);
   ix41524 : inv02 port map ( Y=>nx41525, A=>nx42971);
   ix41526 : inv02 port map ( Y=>nx41527, A=>nx42971);
   ix41528 : inv02 port map ( Y=>nx41529, A=>nx42971);
   ix41530 : buf02 port map ( Y=>nx41531, A=>max_calc_answer_0);
   ix41532 : buf02 port map ( Y=>nx41533, A=>max_calc_answer_0);
   ix41534 : inv02 port map ( Y=>nx41535, A=>nx43137);
   ix41562 : inv02 port map ( Y=>nx41563, A=>nx43155);
   ix41564 : inv02 port map ( Y=>nx41565, A=>nx43031);
   ix41576 : inv02 port map ( Y=>nx41577, A=>nx41575);
   ix41578 : inv02 port map ( Y=>nx41579, A=>nx42975);
   ix41580 : inv02 port map ( Y=>nx41581, A=>nx42975);
   ix41582 : inv02 port map ( Y=>nx41583, A=>nx42975);
   ix41584 : inv02 port map ( Y=>nx41585, A=>nx42975);
   ix41586 : inv02 port map ( Y=>nx41587, A=>nx42539);
   ix41588 : inv02 port map ( Y=>nx41589, A=>nx42539);
   ix41590 : inv02 port map ( Y=>nx41591, A=>nx42539);
   ix41592 : inv02 port map ( Y=>nx41593, A=>nx43205);
   ix41594 : inv02 port map ( Y=>nx41595, A=>nx43205);
   ix41596 : inv02 port map ( Y=>nx41597, A=>nx43205);
   ix41598 : inv02 port map ( Y=>nx41599, A=>nx43205);
   ix41600 : inv02 port map ( Y=>nx41601, A=>nx43205);
   ix41602 : inv02 port map ( Y=>nx41603, A=>nx43205);
   ix41604 : inv02 port map ( Y=>nx41605, A=>nx43205);
   ix41606 : inv02 port map ( Y=>nx41607, A=>nx43209);
   ix41608 : inv02 port map ( Y=>nx41609, A=>nx43209);
   ix41610 : inv02 port map ( Y=>nx41611, A=>nx43209);
   ix41612 : inv02 port map ( Y=>nx41613, A=>nx43209);
   ix41614 : inv02 port map ( Y=>nx41615, A=>nx43209);
   ix41616 : inv02 port map ( Y=>nx41617, A=>nx43209);
   ix41618 : inv02 port map ( Y=>nx41619, A=>nx43209);
   ix41620 : inv02 port map ( Y=>nx41621, A=>nx43213);
   ix41622 : inv02 port map ( Y=>nx41623, A=>nx43213);
   ix41624 : inv02 port map ( Y=>nx41625, A=>nx43213);
   ix41626 : inv02 port map ( Y=>nx41627, A=>nx43213);
   ix41628 : inv02 port map ( Y=>nx41629, A=>nx43213);
   ix41630 : inv02 port map ( Y=>nx41631, A=>nx43213);
   ix41632 : inv02 port map ( Y=>nx41633, A=>nx43213);
   ix41634 : inv02 port map ( Y=>nx41635, A=>nx43217);
   ix41636 : inv02 port map ( Y=>nx41637, A=>nx43217);
   ix41638 : inv02 port map ( Y=>nx41639, A=>nx43217);
   ix41640 : inv02 port map ( Y=>nx41641, A=>nx43217);
   ix41642 : inv02 port map ( Y=>nx41643, A=>nx43217);
   ix41644 : inv02 port map ( Y=>nx41645, A=>nx43217);
   ix41646 : inv02 port map ( Y=>nx41647, A=>nx43217);
   ix41648 : inv02 port map ( Y=>nx41649, A=>nx42549);
   ix41650 : inv02 port map ( Y=>nx41651, A=>nx42549);
   ix41652 : inv02 port map ( Y=>nx41653, A=>nx42549);
   ix41654 : inv02 port map ( Y=>nx41655, A=>nx42549);
   ix41656 : inv02 port map ( Y=>nx41657, A=>nx42549);
   ix41658 : inv02 port map ( Y=>nx41659, A=>nx42549);
   ix41660 : inv02 port map ( Y=>nx41661, A=>nx42443);
   ix41662 : inv02 port map ( Y=>nx41663, A=>nx42445);
   ix41664 : inv02 port map ( Y=>nx41665, A=>nx42445);
   ix41666 : inv02 port map ( Y=>nx41667, A=>nx42445);
   ix41668 : inv02 port map ( Y=>nx41669, A=>nx42445);
   ix41670 : inv02 port map ( Y=>nx41671, A=>nx42445);
   ix41672 : inv02 port map ( Y=>nx41673, A=>nx42445);
   ix41674 : inv02 port map ( Y=>nx41675, A=>nx42445);
   ix41676 : inv02 port map ( Y=>nx41677, A=>nx42447);
   ix41678 : inv02 port map ( Y=>nx41679, A=>nx42447);
   ix41680 : inv02 port map ( Y=>nx41681, A=>nx42447);
   ix41682 : inv02 port map ( Y=>nx41683, A=>nx42447);
   ix41684 : inv02 port map ( Y=>nx41685, A=>nx42447);
   ix41686 : inv02 port map ( Y=>nx41687, A=>nx42447);
   ix41688 : inv02 port map ( Y=>nx41689, A=>nx42447);
   ix41690 : inv02 port map ( Y=>nx41691, A=>nx42449);
   ix41692 : inv02 port map ( Y=>nx41693, A=>nx42449);
   ix41694 : inv02 port map ( Y=>nx41695, A=>nx42449);
   ix41696 : inv02 port map ( Y=>nx41697, A=>nx42449);
   ix41698 : inv02 port map ( Y=>nx41699, A=>nx42449);
   ix41700 : inv02 port map ( Y=>nx41701, A=>nx42449);
   ix41702 : inv02 port map ( Y=>nx41703, A=>nx42449);
   ix41704 : inv02 port map ( Y=>nx41705, A=>nx42451);
   ix41706 : inv02 port map ( Y=>nx41707, A=>nx43123);
   ix41720 : inv02 port map ( Y=>nx41721, A=>nx43131);
   ix41728 : buf02 port map ( Y=>nx41729, A=>neuron_11);
   ix41730 : buf02 port map ( Y=>nx41731, A=>neuron_11);
   ix41740 : buf02 port map ( Y=>nx41741, A=>neuron_10);
   ix41742 : buf02 port map ( Y=>nx41743, A=>neuron_10);
   ix41744 : buf02 port map ( Y=>nx41745, A=>neuron_9);
   ix41746 : buf02 port map ( Y=>nx41747, A=>neuron_9);
   ix41748 : buf02 port map ( Y=>nx41749, A=>neuron_8);
   ix41750 : buf02 port map ( Y=>nx41751, A=>neuron_8);
   ix41752 : buf02 port map ( Y=>nx41753, A=>neuron_7);
   ix41754 : buf02 port map ( Y=>nx41755, A=>neuron_7);
   ix41756 : buf02 port map ( Y=>nx41757, A=>neuron_6);
   ix41758 : buf02 port map ( Y=>nx41759, A=>neuron_6);
   ix41760 : buf02 port map ( Y=>nx41761, A=>neuron_5);
   ix41762 : buf02 port map ( Y=>nx41763, A=>neuron_5);
   ix41764 : buf02 port map ( Y=>nx41765, A=>neuron_4);
   ix41766 : buf02 port map ( Y=>nx41767, A=>neuron_4);
   ix41768 : buf02 port map ( Y=>nx41769, A=>neuron_3);
   ix41770 : buf02 port map ( Y=>nx41771, A=>neuron_3);
   ix41772 : buf02 port map ( Y=>nx41773, A=>neuron_2);
   ix41774 : buf02 port map ( Y=>nx41775, A=>neuron_2);
   ix41776 : buf02 port map ( Y=>nx41777, A=>neuron_1);
   ix41778 : buf02 port map ( Y=>nx41779, A=>neuron_1);
   ix41780 : buf02 port map ( Y=>nx41781, A=>neuron_0);
   ix41782 : buf02 port map ( Y=>nx41783, A=>neuron_0);
   ix41784 : inv02 port map ( Y=>nx41785, A=>nx33026);
   ix41786 : inv02 port map ( Y=>nx41787, A=>nx33026);
   ix41788 : inv01 port map ( Y=>nx41789, A=>nx33023);
   ix41790 : inv01 port map ( Y=>nx41791, A=>nx33023);
   ix41792 : inv01 port map ( Y=>nx41793, A=>nx33023);
   ix41794 : buf02 port map ( Y=>nx41795, A=>neuron_15);
   ix41796 : buf02 port map ( Y=>nx41797, A=>neuron_15);
   ix41798 : buf02 port map ( Y=>nx41799, A=>neuron_14);
   ix41800 : buf02 port map ( Y=>nx41801, A=>neuron_14);
   ix41802 : buf02 port map ( Y=>nx41803, A=>neuron_13);
   ix41804 : buf02 port map ( Y=>nx41805, A=>neuron_13);
   ix41806 : buf02 port map ( Y=>nx41807, A=>neuron_12);
   ix41808 : buf02 port map ( Y=>nx41809, A=>neuron_12);
   ix41810 : inv02 port map ( Y=>nx41811, A=>nx43203);
   ix41812 : inv02 port map ( Y=>nx41813, A=>nx43203);
   ix41814 : inv02 port map ( Y=>nx41815, A=>nx43203);
   ix41816 : inv02 port map ( Y=>nx41817, A=>nx43203);
   ix41818 : inv02 port map ( Y=>nx41819, A=>nx42529);
   ix41832 : inv02 port map ( Y=>nx41833, A=>nx43189);
   ix41846 : inv02 port map ( Y=>nx41847, A=>nx43197);
   ix41854 : inv02 port map ( Y=>nx41855, A=>nx34379);
   ix41856 : inv02 port map ( Y=>nx41857, A=>nx34379);
   ix41858 : inv01 port map ( Y=>nx41859, A=>nx34374);
   ix41860 : inv01 port map ( Y=>nx41861, A=>nx34374);
   ix41862 : inv01 port map ( Y=>nx41863, A=>nx34374);
   ix41864 : inv02 port map ( Y=>nx41865, A=>nx43163);
   ix41878 : inv02 port map ( Y=>nx41879, A=>nx43171);
   ix41886 : inv02 port map ( Y=>nx41887, A=>nx33714);
   ix41888 : inv02 port map ( Y=>nx41889, A=>nx33714);
   ix41890 : inv01 port map ( Y=>nx41891, A=>nx33709);
   ix41892 : inv01 port map ( Y=>nx41893, A=>nx33709);
   ix41894 : inv01 port map ( Y=>nx41895, A=>nx33709);
   ix41904 : inv02 port map ( Y=>nx41905, A=>nx43221);
   ix41918 : inv02 port map ( Y=>nx41919, A=>nx43229);
   ix41926 : inv02 port map ( Y=>nx41927, A=>nx35249);
   ix41928 : inv02 port map ( Y=>nx41929, A=>nx35249);
   ix41930 : inv01 port map ( Y=>nx41931, A=>nx35244);
   ix41932 : inv01 port map ( Y=>nx41933, A=>nx35244);
   ix41934 : inv01 port map ( Y=>nx41935, A=>nx35244);
   ix41936 : inv02 port map ( Y=>nx41937, A=>nx43235);
   ix41950 : inv02 port map ( Y=>nx41951, A=>nx43243);
   ix41958 : inv02 port map ( Y=>nx41959, A=>nx35887);
   ix41960 : inv02 port map ( Y=>nx41961, A=>nx35887);
   ix41962 : inv01 port map ( Y=>nx41963, A=>nx35882);
   ix41964 : inv01 port map ( Y=>nx41965, A=>nx35882);
   ix41966 : inv01 port map ( Y=>nx41967, A=>nx35882);
   ix41968 : inv02 port map ( Y=>nx41969, A=>nx43249);
   ix41982 : inv02 port map ( Y=>nx41983, A=>nx43257);
   ix41990 : inv02 port map ( Y=>nx41991, A=>nx36524);
   ix41992 : inv02 port map ( Y=>nx41993, A=>nx36524);
   ix41994 : inv01 port map ( Y=>nx41995, A=>nx36519);
   ix41996 : inv01 port map ( Y=>nx41997, A=>nx36519);
   ix41998 : inv01 port map ( Y=>nx41999, A=>nx36519);
   ix42000 : inv02 port map ( Y=>nx42001, A=>nx43269);
   ix42014 : inv02 port map ( Y=>nx42015, A=>nx43277);
   ix42022 : inv02 port map ( Y=>nx42023, A=>nx37160);
   ix42024 : inv02 port map ( Y=>nx42025, A=>nx37160);
   ix42026 : inv01 port map ( Y=>nx42027, A=>nx37155);
   ix42028 : inv01 port map ( Y=>nx42029, A=>nx37155);
   ix42030 : inv01 port map ( Y=>nx42031, A=>nx37155);
   ix42040 : inv02 port map ( Y=>nx42041, A=>nx43291);
   ix42054 : inv02 port map ( Y=>nx42055, A=>nx43299);
   ix42062 : inv02 port map ( Y=>nx42063, A=>nx38039);
   ix42064 : inv02 port map ( Y=>nx42065, A=>nx38039);
   ix42066 : inv01 port map ( Y=>nx42067, A=>nx38034);
   ix42068 : inv01 port map ( Y=>nx42069, A=>nx38034);
   ix42070 : inv01 port map ( Y=>nx42071, A=>nx38034);
   ix42072 : inv02 port map ( Y=>nx42073, A=>nx43305);
   ix42086 : inv02 port map ( Y=>nx42087, A=>nx43313);
   ix42094 : inv02 port map ( Y=>nx42095, A=>nx38676);
   ix42096 : inv02 port map ( Y=>nx42097, A=>nx38676);
   ix42098 : inv01 port map ( Y=>nx42099, A=>nx38671);
   ix42100 : inv01 port map ( Y=>nx42101, A=>nx38671);
   ix42102 : inv01 port map ( Y=>nx42103, A=>nx38671);
   ix42104 : inv02 port map ( Y=>nx42105, A=>nx43319);
   ix42118 : inv02 port map ( Y=>nx42119, A=>nx43327);
   ix42126 : inv02 port map ( Y=>nx42127, A=>nx39310);
   ix42128 : inv02 port map ( Y=>nx42129, A=>nx39310);
   ix42130 : inv01 port map ( Y=>nx42131, A=>nx39305);
   ix42132 : inv01 port map ( Y=>nx42133, A=>nx39305);
   ix42134 : inv01 port map ( Y=>nx42135, A=>nx39305);
   ix42160 : buf02 port map ( Y=>nx42161, A=>max_calc_answer_1);
   ix42162 : buf02 port map ( Y=>nx42163, A=>max_calc_answer_1);
   ix42164 : buf02 port map ( Y=>nx42165, A=>max_calc_answer_2);
   ix42166 : buf02 port map ( Y=>nx42167, A=>max_calc_answer_2);
   ix42168 : buf02 port map ( Y=>nx42169, A=>max_calc_answer_3);
   ix42170 : buf02 port map ( Y=>nx42171, A=>max_calc_answer_3);
   ix42172 : buf02 port map ( Y=>nx42173, A=>max_calc_answer_4);
   ix42174 : buf02 port map ( Y=>nx42175, A=>max_calc_answer_4);
   ix42176 : buf02 port map ( Y=>nx42177, A=>max_calc_answer_5);
   ix42178 : buf02 port map ( Y=>nx42179, A=>max_calc_answer_5);
   ix42180 : buf02 port map ( Y=>nx42181, A=>max_calc_answer_6);
   ix42182 : buf02 port map ( Y=>nx42183, A=>max_calc_answer_6);
   ix42184 : buf02 port map ( Y=>nx42185, A=>max_calc_answer_7);
   ix42186 : buf02 port map ( Y=>nx42187, A=>max_calc_answer_7);
   ix42188 : buf02 port map ( Y=>nx42189, A=>max_calc_answer_8);
   ix42190 : buf02 port map ( Y=>nx42191, A=>max_calc_answer_8);
   ix42192 : buf02 port map ( Y=>nx42193, A=>max_calc_answer_9);
   ix42194 : buf02 port map ( Y=>nx42195, A=>max_calc_answer_9);
   ix42196 : buf02 port map ( Y=>nx42197, A=>max_calc_answer_10);
   ix42198 : buf02 port map ( Y=>nx42199, A=>max_calc_answer_10);
   ix42200 : buf02 port map ( Y=>nx42201, A=>max_calc_answer_11);
   ix42202 : buf02 port map ( Y=>nx42203, A=>max_calc_answer_11);
   ix42204 : buf02 port map ( Y=>nx42205, A=>max_calc_answer_12);
   ix42206 : buf02 port map ( Y=>nx42207, A=>max_calc_answer_12);
   ix42208 : buf02 port map ( Y=>nx42209, A=>max_calc_answer_13);
   ix42210 : buf02 port map ( Y=>nx42211, A=>max_calc_answer_13);
   ix42212 : buf02 port map ( Y=>nx42213, A=>max_calc_answer_14);
   ix42214 : buf02 port map ( Y=>nx42215, A=>max_calc_answer_14);
   ix42216 : buf02 port map ( Y=>nx42217, A=>max_calc_answer_15);
   ix42218 : buf02 port map ( Y=>nx42219, A=>max_calc_answer_15);
   ix42226 : inv02 port map ( Y=>nx42227, A=>max_calc_state_2);
   ix42228 : inv02 port map ( Y=>nx42229, A=>nx42803);
   ix42230 : inv02 port map ( Y=>nx42231, A=>nx42803);
   ix42232 : inv02 port map ( Y=>nx42233, A=>nx42803);
   ix42234 : inv02 port map ( Y=>nx42235, A=>nx42803);
   ix42236 : inv02 port map ( Y=>nx42237, A=>nx42803);
   ix42238 : inv02 port map ( Y=>nx42239, A=>nx42803);
   ix42240 : inv02 port map ( Y=>nx42241, A=>nx42803);
   ix42242 : inv02 port map ( Y=>nx42243, A=>nx43389);
   ix42244 : inv02 port map ( Y=>nx42245, A=>nx43389);
   ix42246 : inv02 port map ( Y=>nx42247, A=>nx43389);
   ix42248 : inv02 port map ( Y=>nx42249, A=>nx18145);
   ix42250 : inv02 port map ( Y=>nx42251, A=>nx42847);
   ix42252 : inv02 port map ( Y=>nx42253, A=>nx42847);
   ix42254 : inv02 port map ( Y=>nx42255, A=>nx42847);
   ix42256 : inv02 port map ( Y=>nx42257, A=>nx42847);
   ix42258 : inv02 port map ( Y=>nx42259, A=>sub_state_2);
   ix42260 : inv02 port map ( Y=>nx42261, A=>sub_state_2);
   ix42270 : buf02 port map ( Y=>nx42271, A=>nx31978);
   ix42272 : inv02 port map ( Y=>nx42273, A=>nx18158);
   ix42276 : inv02 port map ( Y=>nx42277, A=>nx4);
   ix42278 : inv02 port map ( Y=>nx42279, A=>nx42855);
   ix42280 : inv02 port map ( Y=>nx42281, A=>nx42855);
   ix42282 : inv02 port map ( Y=>nx42283, A=>nx42855);
   ix42284 : inv02 port map ( Y=>nx42285, A=>enable_decoder_dst_booth);
   ix42286 : inv02 port map ( Y=>nx42287, A=>nx43445);
   ix42288 : inv02 port map ( Y=>nx42289, A=>nx43445);
   ix42290 : inv02 port map ( Y=>nx42291, A=>nx43445);
   ix42292 : inv02 port map ( Y=>nx42293, A=>nx43445);
   ix42294 : inv02 port map ( Y=>nx42295, A=>alu_sel);
   ix42298 : inv02 port map ( Y=>nx42299, A=>nx68);
   ix42300 : inv02 port map ( Y=>nx42301, A=>nx68);
   ix42312 : inv02 port map ( Y=>nx42313, A=>nx42311);
   ix42314 : inv02 port map ( Y=>nx42315, A=>nx43113);
   ix42316 : inv02 port map ( Y=>nx42317, A=>nx43113);
   ix42372 : inv02 port map ( Y=>nx42373, A=>
      booth_booth_integrtaion_0_shift_reg_output_9);
   ix42374 : inv02 port map ( Y=>nx42375, A=>nx43463);
   ix42376 : inv02 port map ( Y=>nx42377, A=>nx43463);
   ix42378 : inv02 port map ( Y=>nx42379, A=>nx43463);
   ix42380 : inv02 port map ( Y=>nx42381, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix42382 : inv02 port map ( Y=>nx42383, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix42384 : buf02 port map ( Y=>nx42385, A=>nx33039);
   ix42386 : buf02 port map ( Y=>nx42387, A=>nx33072);
   ix42388 : buf02 port map ( Y=>nx42389, A=>nx33106);
   ix42390 : buf02 port map ( Y=>nx42391, A=>nx33140);
   ix42392 : buf02 port map ( Y=>nx42393, A=>nx33174);
   ix42394 : buf02 port map ( Y=>nx42395, A=>nx33208);
   ix42396 : buf02 port map ( Y=>nx42397, A=>nx33244);
   ix42442 : inv02 port map ( Y=>nx42443, A=>nx43437);
   ix42444 : inv02 port map ( Y=>nx42445, A=>nx43437);
   ix42446 : inv02 port map ( Y=>nx42447, A=>nx43437);
   ix42448 : inv02 port map ( Y=>nx42449, A=>nx43437);
   ix42450 : inv02 port map ( Y=>nx42451, A=>nx43437);
   ix42452 : inv02 port map ( Y=>nx42453, A=>max_calc_state_1);
   ix42454 : inv02 port map ( Y=>nx42455, A=>nx43453);
   ix42456 : inv02 port map ( Y=>nx42457, A=>nx43453);
   ix42458 : inv02 port map ( Y=>nx42459, A=>
      booth_booth_integrtaion_9_shift_reg_output_9);
   ix42460 : inv02 port map ( Y=>nx42461, A=>nx43471);
   ix42462 : inv02 port map ( Y=>nx42463, A=>nx43471);
   ix42464 : inv02 port map ( Y=>nx42465, A=>nx43471);
   ix42466 : inv02 port map ( Y=>nx42467, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix42468 : inv02 port map ( Y=>nx42469, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix42470 : buf02 port map ( Y=>nx42471, A=>nx33727);
   ix42472 : buf02 port map ( Y=>nx42473, A=>nx33762);
   ix42474 : buf02 port map ( Y=>nx42475, A=>nx33798);
   ix42476 : buf02 port map ( Y=>nx42477, A=>nx33834);
   ix42478 : buf02 port map ( Y=>nx42479, A=>nx33870);
   ix42480 : buf02 port map ( Y=>nx42481, A=>nx33906);
   ix42482 : buf02 port map ( Y=>nx42483, A=>nx33944);
   ix42496 : inv02 port map ( Y=>nx42497, A=>
      booth_booth_integrtaion_8_shift_reg_output_9);
   ix42498 : inv02 port map ( Y=>nx42499, A=>nx43467);
   ix42500 : inv02 port map ( Y=>nx42501, A=>nx43467);
   ix42502 : inv02 port map ( Y=>nx42503, A=>nx43467);
   ix42504 : inv02 port map ( Y=>nx42505, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix42506 : inv02 port map ( Y=>nx42507, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix42508 : buf02 port map ( Y=>nx42509, A=>nx34392);
   ix42510 : buf02 port map ( Y=>nx42511, A=>nx34427);
   ix42512 : buf02 port map ( Y=>nx42513, A=>nx34463);
   ix42514 : buf02 port map ( Y=>nx42515, A=>nx34499);
   ix42516 : buf02 port map ( Y=>nx42517, A=>nx34535);
   ix42518 : buf02 port map ( Y=>nx42519, A=>nx34571);
   ix42520 : buf02 port map ( Y=>nx42521, A=>nx34609);
   ix42526 : inv02 port map ( Y=>nx42527, A=>nx2862);
   ix42528 : inv02 port map ( Y=>nx42529, A=>nx42871);
   ix42538 : inv02 port map ( Y=>nx42539, A=>nx43391);
   ix42540 : inv02 port map ( Y=>nx42541, A=>nx43459);
   ix42542 : inv02 port map ( Y=>nx42543, A=>nx43459);
   ix42544 : inv02 port map ( Y=>nx42545, A=>nx43459);
   ix42546 : inv02 port map ( Y=>nx42547, A=>nx43459);
   ix42548 : inv02 port map ( Y=>nx42549, A=>nx43459);
   ix42550 : inv02 port map ( Y=>nx42551, A=>
      booth_booth_integrtaion_1_shift_reg_output_9);
   ix42552 : inv02 port map ( Y=>nx42553, A=>nx43475);
   ix42554 : inv02 port map ( Y=>nx42555, A=>nx43475);
   ix42556 : inv02 port map ( Y=>nx42557, A=>nx43475);
   ix42558 : inv02 port map ( Y=>nx42559, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix42560 : inv02 port map ( Y=>nx42561, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix42562 : buf02 port map ( Y=>nx42563, A=>nx35262);
   ix42564 : buf02 port map ( Y=>nx42565, A=>nx35297);
   ix42566 : buf02 port map ( Y=>nx42567, A=>nx35333);
   ix42568 : buf02 port map ( Y=>nx42569, A=>nx35369);
   ix42570 : buf02 port map ( Y=>nx42571, A=>nx35405);
   ix42572 : buf02 port map ( Y=>nx42573, A=>nx35441);
   ix42574 : buf02 port map ( Y=>nx42575, A=>nx35479);
   ix42576 : inv02 port map ( Y=>nx42577, A=>
      booth_booth_integrtaion_2_shift_reg_output_9);
   ix42578 : inv02 port map ( Y=>nx42579, A=>nx43479);
   ix42580 : inv02 port map ( Y=>nx42581, A=>nx43479);
   ix42582 : inv02 port map ( Y=>nx42583, A=>nx43479);
   ix42584 : inv02 port map ( Y=>nx42585, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix42586 : inv02 port map ( Y=>nx42587, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix42588 : buf02 port map ( Y=>nx42589, A=>nx35900);
   ix42590 : buf02 port map ( Y=>nx42591, A=>nx35935);
   ix42592 : buf02 port map ( Y=>nx42593, A=>nx35971);
   ix42594 : buf02 port map ( Y=>nx42595, A=>nx36007);
   ix42596 : buf02 port map ( Y=>nx42597, A=>nx36043);
   ix42598 : buf02 port map ( Y=>nx42599, A=>nx36079);
   ix42600 : buf02 port map ( Y=>nx42601, A=>nx36117);
   ix42602 : inv02 port map ( Y=>nx42603, A=>
      booth_booth_integrtaion_4_shift_reg_output_9);
   ix42604 : inv02 port map ( Y=>nx42605, A=>nx43483);
   ix42606 : inv02 port map ( Y=>nx42607, A=>nx43483);
   ix42608 : inv02 port map ( Y=>nx42609, A=>nx43483);
   ix42610 : inv02 port map ( Y=>nx42611, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix42612 : inv02 port map ( Y=>nx42613, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix42614 : buf02 port map ( Y=>nx42615, A=>nx36537);
   ix42616 : buf02 port map ( Y=>nx42617, A=>nx36572);
   ix42618 : buf02 port map ( Y=>nx42619, A=>nx36608);
   ix42620 : buf02 port map ( Y=>nx42621, A=>nx36644);
   ix42622 : buf02 port map ( Y=>nx42623, A=>nx36680);
   ix42624 : buf02 port map ( Y=>nx42625, A=>nx36716);
   ix42626 : buf02 port map ( Y=>nx42627, A=>nx36754);
   ix42630 : inv02 port map ( Y=>nx42631, A=>nx43341);
   ix42632 : inv02 port map ( Y=>nx42633, A=>nx43341);
   ix42634 : inv02 port map ( Y=>nx42635, A=>nx43341);
   ix42636 : inv02 port map ( Y=>nx42637, A=>nx43341);
   ix42638 : inv02 port map ( Y=>nx42639, A=>nx43341);
   ix42640 : inv02 port map ( Y=>nx42641, A=>nx43263);
   ix42642 : inv02 port map ( Y=>nx42643, A=>nx43263);
   ix42644 : inv02 port map ( Y=>nx42645, A=>nx43263);
   ix42646 : inv02 port map ( Y=>nx42647, A=>nx43263);
   ix42650 : inv02 port map ( Y=>nx42651, A=>
      booth_booth_integrtaion_5_shift_reg_output_9);
   ix42652 : inv02 port map ( Y=>nx42653, A=>nx43487);
   ix42654 : inv02 port map ( Y=>nx42655, A=>nx43487);
   ix42656 : inv02 port map ( Y=>nx42657, A=>nx43487);
   ix42658 : inv02 port map ( Y=>nx42659, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix42660 : inv02 port map ( Y=>nx42661, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix42662 : buf02 port map ( Y=>nx42663, A=>nx37173);
   ix42664 : buf02 port map ( Y=>nx42665, A=>nx37208);
   ix42666 : buf02 port map ( Y=>nx42667, A=>nx37244);
   ix42668 : buf02 port map ( Y=>nx42669, A=>nx37280);
   ix42670 : buf02 port map ( Y=>nx42671, A=>nx37316);
   ix42672 : buf02 port map ( Y=>nx42673, A=>nx37352);
   ix42674 : buf02 port map ( Y=>nx42675, A=>nx37390);
   ix42678 : inv02 port map ( Y=>nx42679, A=>nx42677);
   ix42680 : inv02 port map ( Y=>nx42681, A=>nx42677);
   ix42682 : inv02 port map ( Y=>nx42683, A=>nx42677);
   ix42684 : inv02 port map ( Y=>nx42685, A=>nx42677);
   ix42686 : inv02 port map ( Y=>nx42687, A=>nx42677);
   ix42696 : inv02 port map ( Y=>nx42697, A=>
      booth_booth_integrtaion_3_shift_reg_output_9);
   ix42698 : inv02 port map ( Y=>nx42699, A=>nx43491);
   ix42700 : inv02 port map ( Y=>nx42701, A=>nx43491);
   ix42702 : inv02 port map ( Y=>nx42703, A=>nx43491);
   ix42704 : inv02 port map ( Y=>nx42705, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix42706 : inv02 port map ( Y=>nx42707, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix42708 : buf02 port map ( Y=>nx42709, A=>nx38052);
   ix42710 : buf02 port map ( Y=>nx42711, A=>nx38087);
   ix42712 : buf02 port map ( Y=>nx42713, A=>nx38123);
   ix42714 : buf02 port map ( Y=>nx42715, A=>nx38159);
   ix42716 : buf02 port map ( Y=>nx42717, A=>nx38195);
   ix42718 : buf02 port map ( Y=>nx42719, A=>nx38231);
   ix42720 : buf02 port map ( Y=>nx42721, A=>nx38269);
   ix42722 : inv02 port map ( Y=>nx42723, A=>
      booth_booth_integrtaion_6_shift_reg_output_9);
   ix42724 : inv02 port map ( Y=>nx42725, A=>nx43495);
   ix42726 : inv02 port map ( Y=>nx42727, A=>nx43495);
   ix42728 : inv02 port map ( Y=>nx42729, A=>nx43495);
   ix42730 : inv02 port map ( Y=>nx42731, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix42732 : inv02 port map ( Y=>nx42733, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix42734 : buf02 port map ( Y=>nx42735, A=>nx38689);
   ix42736 : buf02 port map ( Y=>nx42737, A=>nx38724);
   ix42738 : buf02 port map ( Y=>nx42739, A=>nx38760);
   ix42740 : buf02 port map ( Y=>nx42741, A=>nx38796);
   ix42742 : buf02 port map ( Y=>nx42743, A=>nx38832);
   ix42744 : buf02 port map ( Y=>nx42745, A=>nx38868);
   ix42746 : buf02 port map ( Y=>nx42747, A=>nx38906);
   ix42748 : inv02 port map ( Y=>nx42749, A=>
      booth_booth_integrtaion_7_shift_reg_output_9);
   ix42750 : inv02 port map ( Y=>nx42751, A=>nx43499);
   ix42752 : inv02 port map ( Y=>nx42753, A=>nx43499);
   ix42754 : inv02 port map ( Y=>nx42755, A=>nx43499);
   ix42756 : inv02 port map ( Y=>nx42757, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix42758 : inv02 port map ( Y=>nx42759, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix42760 : buf02 port map ( Y=>nx42761, A=>nx39323);
   ix42762 : buf02 port map ( Y=>nx42763, A=>nx39358);
   ix42764 : buf02 port map ( Y=>nx42765, A=>nx39394);
   ix42766 : buf02 port map ( Y=>nx42767, A=>nx39430);
   ix42768 : buf02 port map ( Y=>nx42769, A=>nx39466);
   ix42770 : buf02 port map ( Y=>nx42771, A=>nx39502);
   ix42772 : buf02 port map ( Y=>nx42773, A=>nx39540);
   ix42788 : inv02 port map ( Y=>nx42789, A=>nx41469);
   ix42790 : inv02 port map ( Y=>nx42791, A=>nx41469);
   ix42792 : inv02 port map ( Y=>nx42793, A=>nx41469);
   ix42794 : inv02 port map ( Y=>nx42795, A=>nx32729);
   ix42796 : inv02 port map ( Y=>nx42797, A=>nx43503);
   ix42798 : inv02 port map ( Y=>nx42799, A=>nx43503);
   ix42800 : inv02 port map ( Y=>nx42801, A=>nx43503);
   ix42802 : inv02 port map ( Y=>nx42803, A=>nx42227);
   ix42804 : inv02 port map ( Y=>nx42805, A=>nx42227);
   ix42808 : inv02 port map ( Y=>nx42809, A=>nx33312);
   ix42810 : inv02 port map ( Y=>nx42811, A=>nx43511);
   ix42812 : inv02 port map ( Y=>nx42813, A=>nx43511);
   ix42814 : inv02 port map ( Y=>nx42815, A=>nx43511);
   ix42816 : inv02 port map ( Y=>nx42817, A=>ready_signal);
   ix42818 : inv02 port map ( Y=>nx42819, A=>max_calc_state_2);
   ix20935 : or02 port map ( Y=>nx18189, A0=>nx43389, A1=>nx42925);
   ix1701 : or02 port map ( Y=>nx31926, A0=>nx42257, A1=>nx31938);
   ix1659 : and02 port map ( Y=>nx18153, A0=>nx42877, A1=>nx42883);
   ix1657 : and03 port map ( Y=>nx18159, A0=>state_0, A1=>nx42879, A2=>
      nx42883);
   ix19102 : mux21_ni port map ( Y=>nx19101, A0=>num_in_2, A1=>num_out_2, S0
      =>nx42907);
   ix19092 : mux21_ni port map ( Y=>nx19091, A0=>num_in_2, A1=>nx570, S0=>
      nx43107);
   ix571 : ao22 port map ( Y=>nx570, A0=>data_in(2), A1=>nx68, B0=>nx18162, 
      B1=>nx42855);
   ix18872 : mux21 port map ( Y=>nx18871, A0=>nx43097, A1=>nx42283, S0=>
      nx43049);
   ix31954 : and03 port map ( Y=>nx42263, A0=>nx31955, A1=>nx31957, A2=>
      nx246);
   ix31962 : and03 port map ( Y=>nx31961, A0=>nx42887, A1=>nx43041, A2=>
      nx42891);
   ix31967 : xnor2 port map ( Y=>nx31966, A0=>nx42891, A1=>nx42887);
   ix31975 : and03 port map ( Y=>nx31974, A0=>nx42887, A1=>nx43041, A2=>
      nx42861);
   ix1583 : and02 port map ( Y=>nx1582, A0=>nx42847, A1=>nx42867);
   ix31982 : nand02 port map ( Y=>nx18158, A0=>nx42897, A1=>nx42789);
   ix18662 : mux21 port map ( Y=>nx18661, A0=>nx42283, A1=>nx41469, S0=>
      nx31991);
   ix133 : mux21 port map ( Y=>nx132, A0=>nx122, A1=>nx42277, S0=>nx42257);
   ix31995 : nor03_2x port map ( Y=>nx4, A0=>nx31906, A1=>state_2, A2=>
      nx42885);
   ix18852 : mux21_ni port map ( Y=>nx18851, A0=>nx41421, A1=>output_17, S0
      =>nx42897);
   ix18842 : mux21_ni port map ( Y=>nx18841, A0=>output_17, A1=>output_16, 
      S0=>nx42897);
   ix18832 : mux21_ni port map ( Y=>nx18831, A0=>output_16, A1=>output_15, 
      S0=>nx42897);
   ix18822 : mux21_ni port map ( Y=>nx18821, A0=>output_15, A1=>output_14, 
      S0=>nx42899);
   ix18812 : mux21_ni port map ( Y=>nx18811, A0=>output_14, A1=>output_13, 
      S0=>nx42899);
   ix18802 : mux21_ni port map ( Y=>nx18801, A0=>output_13, A1=>output_12, 
      S0=>nx42899);
   ix18792 : mux21_ni port map ( Y=>nx18791, A0=>output_12, A1=>output_11, 
      S0=>nx42899);
   ix18782 : mux21_ni port map ( Y=>nx18781, A0=>output_11, A1=>output_10, 
      S0=>nx42899);
   ix18772 : mux21_ni port map ( Y=>nx18771, A0=>output_10, A1=>output_9, S0
      =>nx42899);
   ix18762 : mux21_ni port map ( Y=>nx18761, A0=>output_9, A1=>output_8, S0
      =>nx42899);
   ix18752 : mux21_ni port map ( Y=>nx18751, A0=>output_8, A1=>output_7, S0
      =>nx42901);
   ix18742 : mux21_ni port map ( Y=>nx18741, A0=>output_7, A1=>output_6, S0
      =>nx42901);
   ix18732 : mux21_ni port map ( Y=>nx18731, A0=>output_6, A1=>output_5, S0
      =>nx42901);
   ix18722 : mux21_ni port map ( Y=>nx18721, A0=>output_5, A1=>output_4, S0
      =>nx42901);
   ix18712 : mux21_ni port map ( Y=>nx18711, A0=>output_4, A1=>output_3, S0
      =>nx42901);
   ix18702 : mux21_ni port map ( Y=>nx18701, A0=>output_3, A1=>output_2, S0
      =>nx42901);
   ix18692 : mux21_ni port map ( Y=>nx18691, A0=>output_2, A1=>output_1, S0
      =>nx42901);
   ix18682 : mux21_ni port map ( Y=>nx18681, A0=>output_1, A1=>output_0, S0
      =>nx42903);
   ix1665 : ao21 port map ( Y=>nx18146, A0=>nx31906, A1=>nx42885, B0=>
      nx42879);
   ix1643 : and03 port map ( Y=>nx18155, A0=>nx31906, A1=>state_2, A2=>
      nx42885);
   ix37 : or03 port map ( Y=>nx36, A0=>nx42889, A1=>sub_state_2, A2=>nx42861
   );
   ix19032 : mux21_ni port map ( Y=>nx19031, A0=>alu_inp1_1, A1=>nx500, S0=>
      nx43049);
   ix501 : mux21_ni port map ( Y=>nx500, A0=>address_out(1), A1=>num_out_1, 
      S0=>nx42855);
   ix19022 : mux21_ni port map ( Y=>nx19021, A0=>num_in_1, A1=>num_out_1, S0
      =>nx42907);
   ix19012 : mux21 port map ( Y=>nx19011, A0=>nx32150, A1=>nx32072, S0=>
      nx43107);
   ix69 : and03 port map ( Y=>nx68, A0=>nx31906, A1=>nx42879, A2=>nx42885);
   ix443 : mux21_ni port map ( Y=>nx442, A0=>alu_inp1_0, A1=>nx41413, S0=>
      nx32089);
   ix18952 : mux21_ni port map ( Y=>nx18951, A0=>alu_inp1_0, A1=>nx420, S0=>
      nx43049);
   ix421 : mux21_ni port map ( Y=>nx420, A0=>address_out(0), A1=>num_out_0, 
      S0=>nx42855);
   ix18942 : mux21_ni port map ( Y=>nx18941, A0=>num_in_0, A1=>num_out_0, S0
      =>nx42907);
   ix18932 : mux21_ni port map ( Y=>nx18931, A0=>num_in_0, A1=>nx406, S0=>
      nx43107);
   ix407 : ao22 port map ( Y=>nx406, A0=>data_in(0), A1=>nx68, B0=>nx360, B1
      =>nx42855);
   ix32086 : xor2 port map ( Y=>nx32085, A0=>alu_inp1_0, A1=>nx32089);
   ix18962 : or02 port map ( Y=>nx18961, A0=>alu_inp2_0, A1=>nx43049);
   ix32096 : and03 port map ( Y=>nx42303, A0=>nx86, A1=>nx31955, A2=>nx31959
   );
   ix87 : mux21 port map ( Y=>nx86, A0=>nx43041, A1=>nx42283, S0=>nx42301);
   ix18922 : mux21_ni port map ( Y=>nx18921, A0=>address_in_0, A1=>
      address_out(0), S0=>nx42915);
   ix18912 : mux21_ni port map ( Y=>nx18911, A0=>address_in_0, A1=>nx388, S0
      =>nx43117);
   ix32112 : oai21 port map ( Y=>nx42311, A0=>nx42889, A1=>nx42301, B0=>
      nx33299);
   ix32114 : mux21 port map ( Y=>nx32113, A0=>temp_0, A1=>neuron_address_0, 
      S0=>nx43043);
   ix18892 : mux21_ni port map ( Y=>nx18891, A0=>nx362, A1=>neuron_address_0, 
      S0=>nx42971);
   ix363 : nor02ii port map ( Y=>nx362, A0=>nx32085, A1=>nx42847);
   ix359 : nand04 port map ( Y=>nx41521, A0=>nx42847, A1=>nx42825, A2=>
      nx42867, A3=>nx42881);
   ix42824 : inv01 port map ( Y=>nx42825, A=>nx32119);
   ix32120 : or03 port map ( Y=>nx32119, A0=>nx42891, A1=>sub_state_2, A2=>
      nx42889);
   ix18902 : mux21_ni port map ( Y=>nx18901, A0=>nx360, A1=>temp_0, S0=>
      nx42965);
   ix285 : and03 port map ( Y=>nx284, A0=>nx31966, A1=>nx42867, A2=>nx42881
   );
   ix337 : and03 port map ( Y=>nx336, A0=>nx42879, A1=>nx42885, A2=>nx31906
   );
   ix307 : and02 port map ( Y=>nx306, A0=>nx42867, A1=>nx42881);
   ix32149 : xor2 port map ( Y=>nx32148, A0=>alu_inp1_1, A1=>nx43097);
   ix19002 : mux21_ni port map ( Y=>nx19001, A0=>address_in_1, A1=>
      address_out(1), S0=>nx42915);
   ix18992 : mux21_ni port map ( Y=>nx18991, A0=>address_in_1, A1=>nx468, S0
      =>nx43117);
   ix469 : ao22 port map ( Y=>nx468, A0=>nx444, A1=>nx43113, B0=>nx42849, B1
      =>nx42827);
   ix32161 : mux21_ni port map ( Y=>nx42827, A0=>temp_1, A1=>
      neuron_address_1, S0=>nx43043);
   ix18982 : mux21_ni port map ( Y=>nx18981, A0=>nx444, A1=>temp_1, S0=>
      nx42965);
   ix32176 : xnor2 port map ( Y=>nx32175, A0=>nx32197, A1=>nx43097);
   ix19082 : mux21_ni port map ( Y=>nx19081, A0=>alu_inp1_2, A1=>nx554, S0=>
      nx43049);
   ix555 : mux21_ni port map ( Y=>nx554, A0=>address_out(2), A1=>num_out_2, 
      S0=>nx42857);
   ix19072 : mux21_ni port map ( Y=>nx19071, A0=>address_in_2, A1=>
      address_out(2), S0=>nx42915);
   ix19062 : mux21_ni port map ( Y=>nx19061, A0=>address_in_2, A1=>nx538, S0
      =>nx43117);
   ix32186 : mux21 port map ( Y=>nx32185, A0=>temp_2, A1=>neuron_address_2, 
      S0=>nx43043);
   ix19042 : mux21_ni port map ( Y=>nx19041, A0=>nx516, A1=>neuron_address_2, 
      S0=>nx42971);
   ix517 : nor02ii port map ( Y=>nx516, A0=>nx31946, A1=>nx42849);
   ix19052 : mux21_ni port map ( Y=>nx19051, A0=>nx18162, A1=>temp_2, S0=>
      nx42965);
   ix19172 : mux21_ni port map ( Y=>nx19171, A0=>num_in_3, A1=>num_out_3, S0
      =>nx42907);
   ix19162 : mux21 port map ( Y=>nx19161, A0=>nx32238, A1=>nx32208, S0=>
      nx43107);
   ix32213 : xor2 port map ( Y=>nx32212, A0=>alu_inp1_3, A1=>nx43099);
   ix19152 : mux21_ni port map ( Y=>nx19151, A0=>alu_inp1_3, A1=>nx636, S0=>
      nx43049);
   ix637 : mux21_ni port map ( Y=>nx636, A0=>address_out(3), A1=>num_out_3, 
      S0=>nx42857);
   ix19142 : mux21_ni port map ( Y=>nx19141, A0=>address_in_3, A1=>
      address_out(3), S0=>nx42915);
   ix19132 : mux21_ni port map ( Y=>nx19131, A0=>address_in_3, A1=>nx620, S0
      =>nx43117);
   ix621 : ao22 port map ( Y=>nx620, A0=>nx18163, A1=>nx43113, B0=>nx42849, 
      B1=>nx42829);
   ix32225 : mux21_ni port map ( Y=>nx42829, A0=>temp_3, A1=>
      neuron_address_3, S0=>nx43043);
   ix19122 : mux21_ni port map ( Y=>nx19121, A0=>nx18163, A1=>temp_3, S0=>
      nx42965);
   ix19242 : mux21_ni port map ( Y=>nx19241, A0=>num_in_4, A1=>num_out_4, S0
      =>nx42907);
   ix19232 : mux21_ni port map ( Y=>nx19231, A0=>num_in_4, A1=>nx724, S0=>
      nx43107);
   ix32252 : xnor2 port map ( Y=>nx32251, A0=>nx32273, A1=>nx43099);
   ix19222 : mux21_ni port map ( Y=>nx19221, A0=>alu_inp1_4, A1=>nx708, S0=>
      nx43049);
   ix709 : mux21_ni port map ( Y=>nx708, A0=>address_out(4), A1=>num_out_4, 
      S0=>nx42857);
   ix19212 : mux21_ni port map ( Y=>nx19211, A0=>address_in_4, A1=>
      address_out(4), S0=>nx42915);
   ix19202 : mux21_ni port map ( Y=>nx19201, A0=>address_in_4, A1=>nx692, S0
      =>nx43117);
   ix32262 : mux21 port map ( Y=>nx32261, A0=>temp_4, A1=>neuron_address_4, 
      S0=>nx43043);
   ix19182 : mux21_ni port map ( Y=>nx19181, A0=>nx670, A1=>neuron_address_4, 
      S0=>nx42971);
   ix671 : nor02ii port map ( Y=>nx670, A0=>nx32246, A1=>nx42849);
   ix19192 : mux21_ni port map ( Y=>nx19191, A0=>nx18165, A1=>temp_4, S0=>
      nx42965);
   ix19312 : mux21_ni port map ( Y=>nx19311, A0=>num_in_5, A1=>num_out_5, S0
      =>nx42907);
   ix19302 : mux21 port map ( Y=>nx19301, A0=>nx32313, A1=>nx32283, S0=>
      nx43107);
   ix32288 : xor2 port map ( Y=>nx32287, A0=>alu_inp1_5, A1=>nx43099);
   ix19292 : mux21_ni port map ( Y=>nx19291, A0=>alu_inp1_5, A1=>nx788, S0=>
      nx43051);
   ix789 : mux21_ni port map ( Y=>nx788, A0=>address_out(5), A1=>num_out_5, 
      S0=>nx42857);
   ix19282 : mux21_ni port map ( Y=>nx19281, A0=>address_in_5, A1=>
      address_out(5), S0=>nx42915);
   ix19272 : mux21_ni port map ( Y=>nx19271, A0=>address_in_5, A1=>nx772, S0
      =>nx43117);
   ix773 : ao22 port map ( Y=>nx772, A0=>nx18167, A1=>nx43113, B0=>nx42849, 
      B1=>nx42831);
   ix32300 : mux21_ni port map ( Y=>nx42831, A0=>temp_5, A1=>
      neuron_address_5, S0=>nx43043);
   ix19262 : mux21_ni port map ( Y=>nx19261, A0=>nx18167, A1=>temp_5, S0=>
      nx42965);
   ix19382 : mux21_ni port map ( Y=>nx19381, A0=>num_in_6, A1=>num_out_6, S0
      =>nx42909);
   ix19372 : mux21_ni port map ( Y=>nx19371, A0=>num_in_6, A1=>nx876, S0=>
      nx43107);
   ix32327 : xnor2 port map ( Y=>nx32326, A0=>nx32348, A1=>nx43099);
   ix19362 : mux21_ni port map ( Y=>nx19361, A0=>alu_inp1_6, A1=>nx860, S0=>
      nx43051);
   ix861 : mux21_ni port map ( Y=>nx860, A0=>address_out(6), A1=>num_out_6, 
      S0=>nx42857);
   ix19352 : mux21_ni port map ( Y=>nx19351, A0=>address_in_6, A1=>
      address_out(6), S0=>nx42917);
   ix19342 : mux21_ni port map ( Y=>nx19341, A0=>address_in_6, A1=>nx844, S0
      =>nx43117);
   ix32337 : mux21 port map ( Y=>nx32336, A0=>temp_6, A1=>neuron_address_6, 
      S0=>nx43043);
   ix19322 : mux21_ni port map ( Y=>nx19321, A0=>nx822, A1=>neuron_address_6, 
      S0=>nx42971);
   ix823 : nor02ii port map ( Y=>nx822, A0=>nx32321, A1=>nx42849);
   ix19332 : mux21_ni port map ( Y=>nx19331, A0=>nx18169, A1=>temp_6, S0=>
      nx42967);
   ix19452 : mux21_ni port map ( Y=>nx19451, A0=>num_in_7, A1=>num_out_7, S0
      =>nx42909);
   ix19442 : mux21 port map ( Y=>nx19441, A0=>nx32387, A1=>nx32357, S0=>
      nx43109);
   ix32362 : xor2 port map ( Y=>nx32361, A0=>alu_inp1_7, A1=>nx43099);
   ix19432 : mux21_ni port map ( Y=>nx19431, A0=>alu_inp1_7, A1=>nx938, S0=>
      nx43051);
   ix939 : mux21_ni port map ( Y=>nx938, A0=>address_out(7), A1=>num_out_7, 
      S0=>nx42857);
   ix19422 : mux21_ni port map ( Y=>nx19421, A0=>address_in_7, A1=>
      address_out(7), S0=>nx42917);
   ix19412 : mux21_ni port map ( Y=>nx19411, A0=>address_in_7, A1=>nx922, S0
      =>nx43119);
   ix923 : ao22 port map ( Y=>nx922, A0=>nx18171, A1=>nx43113, B0=>nx42849, 
      B1=>nx42833);
   ix32374 : mux21_ni port map ( Y=>nx42833, A0=>temp_7, A1=>
      neuron_address_7, S0=>nx43045);
   ix19402 : mux21_ni port map ( Y=>nx19401, A0=>nx18171, A1=>temp_7, S0=>
      nx42967);
   ix19522 : mux21_ni port map ( Y=>nx19521, A0=>num_in_8, A1=>num_out_8, S0
      =>nx42909);
   ix19512 : mux21_ni port map ( Y=>nx19511, A0=>num_in_8, A1=>nx1026, S0=>
      nx43109);
   ix32401 : xnor2 port map ( Y=>nx32400, A0=>nx32422, A1=>nx43099);
   ix19502 : mux21_ni port map ( Y=>nx19501, A0=>alu_inp1_8, A1=>nx1010, S0
      =>nx43051);
   ix1011 : mux21_ni port map ( Y=>nx1010, A0=>address_out(8), A1=>num_out_8, 
      S0=>nx42857);
   ix19492 : mux21_ni port map ( Y=>nx19491, A0=>address_in_8, A1=>
      address_out(8), S0=>nx42917);
   ix19482 : mux21_ni port map ( Y=>nx19481, A0=>address_in_8, A1=>nx994, S0
      =>nx43119);
   ix32411 : mux21 port map ( Y=>nx32410, A0=>temp_8, A1=>neuron_address_8, 
      S0=>nx43045);
   ix19462 : mux21_ni port map ( Y=>nx19461, A0=>nx972, A1=>neuron_address_8, 
      S0=>nx42973);
   ix973 : nor02ii port map ( Y=>nx972, A0=>nx32395, A1=>nx42851);
   ix19472 : mux21_ni port map ( Y=>nx19471, A0=>nx18173, A1=>temp_8, S0=>
      nx42967);
   ix19592 : mux21_ni port map ( Y=>nx19591, A0=>num_in_9, A1=>num_out_9, S0
      =>nx42909);
   ix19582 : mux21 port map ( Y=>nx19581, A0=>nx32462, A1=>nx32432, S0=>
      nx43109);
   ix32437 : xor2 port map ( Y=>nx32436, A0=>alu_inp1_9, A1=>nx43099);
   ix19572 : mux21_ni port map ( Y=>nx19571, A0=>alu_inp1_9, A1=>nx1092, S0
      =>nx43051);
   ix1093 : mux21_ni port map ( Y=>nx1092, A0=>address_out(9), A1=>num_out_9, 
      S0=>nx42859);
   ix19562 : mux21_ni port map ( Y=>nx19561, A0=>address_in_9, A1=>
      address_out(9), S0=>nx42917);
   ix19552 : mux21_ni port map ( Y=>nx19551, A0=>address_in_9, A1=>nx1076, 
      S0=>nx43119);
   ix1077 : ao22 port map ( Y=>nx1076, A0=>nx18175, A1=>nx43113, B0=>nx42851, 
      B1=>nx42835);
   ix32449 : mux21_ni port map ( Y=>nx42835, A0=>temp_9, A1=>
      neuron_address_9, S0=>nx43045);
   ix19542 : mux21_ni port map ( Y=>nx19541, A0=>nx18175, A1=>temp_9, S0=>
      nx42967);
   ix19662 : mux21_ni port map ( Y=>nx19661, A0=>num_in_10, A1=>num_out_10, 
      S0=>nx42909);
   ix19652 : mux21_ni port map ( Y=>nx19651, A0=>num_in_10, A1=>nx1180, S0=>
      nx43109);
   ix32476 : xnor2 port map ( Y=>nx32475, A0=>nx32497, A1=>nx43101);
   ix19642 : mux21_ni port map ( Y=>nx19641, A0=>alu_inp1_10, A1=>nx1164, S0
      =>nx43051);
   ix1165 : mux21_ni port map ( Y=>nx1164, A0=>address_out(10), A1=>
      num_out_10, S0=>nx42859);
   ix19632 : mux21_ni port map ( Y=>nx19631, A0=>address_in_10, A1=>
      address_out(10), S0=>nx42917);
   ix19622 : mux21_ni port map ( Y=>nx19621, A0=>address_in_10, A1=>nx1148, 
      S0=>nx43119);
   ix32486 : mux21 port map ( Y=>nx32485, A0=>temp_10, A1=>neuron_address_10, 
      S0=>nx43045);
   ix19602 : mux21_ni port map ( Y=>nx19601, A0=>nx1126, A1=>
      neuron_address_10, S0=>nx42973);
   ix1127 : nor02ii port map ( Y=>nx1126, A0=>nx32470, A1=>nx42851);
   ix19612 : mux21_ni port map ( Y=>nx19611, A0=>nx18177, A1=>temp_10, S0=>
      nx42967);
   ix19732 : mux21_ni port map ( Y=>nx19731, A0=>num_in_11, A1=>num_out_11, 
      S0=>nx42909);
   ix19722 : mux21 port map ( Y=>nx19721, A0=>nx32536, A1=>nx32506, S0=>
      nx43109);
   ix32511 : xor2 port map ( Y=>nx32510, A0=>alu_inp1_11, A1=>nx43101);
   ix19712 : mux21_ni port map ( Y=>nx19711, A0=>alu_inp1_11, A1=>nx1242, S0
      =>nx43051);
   ix1243 : mux21_ni port map ( Y=>nx1242, A0=>address_out(11), A1=>
      num_out_11, S0=>nx42859);
   ix19702 : mux21_ni port map ( Y=>nx19701, A0=>address_in_11, A1=>
      address_out(11), S0=>nx42917);
   ix19692 : mux21_ni port map ( Y=>nx19691, A0=>address_in_11, A1=>nx1226, 
      S0=>nx43119);
   ix1227 : ao22 port map ( Y=>nx1226, A0=>nx18178, A1=>nx43115, B0=>nx42851, 
      B1=>nx42837);
   ix32523 : mux21_ni port map ( Y=>nx42837, A0=>temp_11, A1=>
      neuron_address_11, S0=>nx43045);
   ix19682 : mux21_ni port map ( Y=>nx19681, A0=>nx18178, A1=>temp_11, S0=>
      nx42967);
   ix19802 : mux21_ni port map ( Y=>nx19801, A0=>num_in_12, A1=>num_out_12, 
      S0=>nx42909);
   ix19792 : mux21_ni port map ( Y=>nx19791, A0=>num_in_12, A1=>nx1330, S0=>
      nx43109);
   ix32550 : xnor2 port map ( Y=>nx32549, A0=>nx32571, A1=>nx43101);
   ix19782 : mux21_ni port map ( Y=>nx19781, A0=>alu_inp1_12, A1=>nx1314, S0
      =>nx43053);
   ix1315 : mux21_ni port map ( Y=>nx1314, A0=>address_out(12), A1=>
      num_out_12, S0=>nx42859);
   ix19772 : mux21_ni port map ( Y=>nx19771, A0=>address_in_12, A1=>
      address_out(12), S0=>nx42917);
   ix19762 : mux21_ni port map ( Y=>nx19761, A0=>address_in_12, A1=>nx1298, 
      S0=>nx43119);
   ix32560 : mux21 port map ( Y=>nx32559, A0=>temp_12, A1=>neuron_address_12, 
      S0=>nx43045);
   ix19742 : mux21_ni port map ( Y=>nx19741, A0=>nx1276, A1=>
      neuron_address_12, S0=>nx42973);
   ix1277 : nor02ii port map ( Y=>nx1276, A0=>nx32544, A1=>nx42851);
   ix19752 : mux21_ni port map ( Y=>nx19751, A0=>nx18179, A1=>temp_12, S0=>
      nx42967);
   ix19872 : mux21_ni port map ( Y=>nx19871, A0=>num_in_13, A1=>num_out_13, 
      S0=>nx42911);
   ix19862 : mux21 port map ( Y=>nx19861, A0=>nx32611, A1=>nx32581, S0=>
      nx43109);
   ix32586 : xor2 port map ( Y=>nx32585, A0=>alu_inp1_13, A1=>nx43101);
   ix19852 : mux21_ni port map ( Y=>nx19851, A0=>alu_inp1_13, A1=>nx1394, S0
      =>nx43053);
   ix1395 : mux21_ni port map ( Y=>nx1394, A0=>address_out(13), A1=>
      num_out_13, S0=>nx42859);
   ix19842 : mux21_ni port map ( Y=>nx19841, A0=>address_in_13, A1=>
      address_out(13), S0=>nx42919);
   ix19832 : mux21_ni port map ( Y=>nx19831, A0=>address_in_13, A1=>nx1378, 
      S0=>nx43119);
   ix1379 : ao22 port map ( Y=>nx1378, A0=>nx18180, A1=>nx43115, B0=>nx42851, 
      B1=>nx42839);
   ix32598 : mux21_ni port map ( Y=>nx42839, A0=>temp_13, A1=>
      neuron_address_13, S0=>nx43045);
   ix19822 : mux21_ni port map ( Y=>nx19821, A0=>nx18180, A1=>temp_13, S0=>
      nx42969);
   ix19942 : mux21_ni port map ( Y=>nx19941, A0=>num_in_14, A1=>num_out_14, 
      S0=>nx42911);
   ix19932 : mux21_ni port map ( Y=>nx19931, A0=>num_in_14, A1=>nx1482, S0=>
      nx43111);
   ix32625 : xnor2 port map ( Y=>nx32624, A0=>nx32646, A1=>nx43101);
   ix19922 : mux21_ni port map ( Y=>nx19921, A0=>alu_inp1_14, A1=>nx1466, S0
      =>nx43053);
   ix1467 : mux21_ni port map ( Y=>nx1466, A0=>address_out(14), A1=>
      num_out_14, S0=>nx42859);
   ix19912 : mux21_ni port map ( Y=>nx19911, A0=>address_in_14, A1=>
      address_out(14), S0=>nx42919);
   ix19902 : mux21_ni port map ( Y=>nx19901, A0=>address_in_14, A1=>nx1450, 
      S0=>nx43121);
   ix32635 : mux21 port map ( Y=>nx32634, A0=>temp_14, A1=>neuron_address_14, 
      S0=>nx42261);
   ix19882 : mux21_ni port map ( Y=>nx19881, A0=>nx1428, A1=>
      neuron_address_14, S0=>nx42973);
   ix1429 : nor02ii port map ( Y=>nx1428, A0=>nx32619, A1=>nx42851);
   ix19892 : mux21_ni port map ( Y=>nx19891, A0=>nx18181, A1=>temp_14, S0=>
      nx42969);
   ix20012 : mux21_ni port map ( Y=>nx20011, A0=>num_in_15, A1=>num_out_15, 
      S0=>nx42911);
   ix20002 : mux21 port map ( Y=>nx20001, A0=>nx32686, A1=>nx32655, S0=>
      nx43111);
   ix32660 : xor2 port map ( Y=>nx32659, A0=>alu_inp1_15, A1=>nx43101);
   ix19992 : mux21_ni port map ( Y=>nx19991, A0=>alu_inp1_15, A1=>nx1544, S0
      =>nx43053);
   ix1545 : mux21_ni port map ( Y=>nx1544, A0=>address_out(15), A1=>
      num_out_15, S0=>nx42859);
   ix19982 : mux21_ni port map ( Y=>nx19981, A0=>address_in_15, A1=>
      address_out(15), S0=>nx42919);
   ix19972 : mux21_ni port map ( Y=>nx19971, A0=>address_in_15, A1=>nx1528, 
      S0=>nx43121);
   ix1529 : ao22 port map ( Y=>nx1528, A0=>nx18182, A1=>nx43115, B0=>nx42853, 
      B1=>nx42841);
   ix32673 : mux21_ni port map ( Y=>nx42841, A0=>temp_15, A1=>
      neuron_address_15, S0=>nx42261);
   ix19962 : mux21_ni port map ( Y=>nx19961, A0=>nx18182, A1=>temp_15, S0=>
      nx42969);
   ix1673 : and02 port map ( Y=>nx1672, A0=>nx42867, A1=>nx31938);
   ix32715 : xor2 port map ( Y=>nx32714, A0=>nx42217, A1=>nx39926);
   ix31812 : mux21_ni port map ( Y=>nx31811, A0=>nx42217, A1=>nx18623, S0=>
      nx43335);
   ix20081 : mux21_ni port map ( Y=>nx18623, A0=>
      max_calc_comparator_first_inp2_15, A1=>
      max_calc_comparator_first_inp1_15, S0=>nx43025);
   ix31622 : mux21_ni port map ( Y=>nx31621, A0=>
      max_calc_comparator_first_inp1_15, A1=>nx20066, S0=>nx43391);
   ix20067 : mux21_ni port map ( Y=>nx20066, A0=>nx20062, A1=>nx20030, S0=>
      nx43031);
   ix20031 : mux21_ni port map ( Y=>nx20030, A0=>max_calc_ans1_15, A1=>
      label_1_output_15, S0=>nx43155);
   ix31582 : mux21_ni port map ( Y=>nx31581, A0=>label_1_output_15, A1=>
      label_1_input_15, S0=>nx43401);
   ix20007 : mux21_ni port map ( Y=>nx20006, A0=>nx20002, A1=>
      label_1_input_state_machine_15, S0=>nx43055);
   ix31572 : mux21_ni port map ( Y=>nx31571, A0=>
      label_1_input_state_machine_15, A1=>data_in(15), S0=>nx43349);
   ix30382 : mux21_ni port map ( Y=>nx30381, A0=>label_1_output_14, A1=>
      label_1_input_14, S0=>nx43401);
   ix18059 : mux21_ni port map ( Y=>nx18058, A0=>nx18054, A1=>
      label_1_input_state_machine_14, S0=>nx43057);
   ix30112 : mux21_ni port map ( Y=>nx30111, A0=>
      label_1_input_state_machine_14, A1=>data_in(14), S0=>nx43349);
   ix30352 : mux21_ni port map ( Y=>nx30351, A0=>label_1_output_12, A1=>
      label_1_input_12, S0=>nx43401);
   ix18001 : mux21_ni port map ( Y=>nx18000, A0=>nx17996, A1=>
      label_1_input_state_machine_12, S0=>nx43057);
   ix30342 : mux21_ni port map ( Y=>nx30341, A0=>
      label_1_input_state_machine_12, A1=>data_in(12), S0=>nx43349);
   ix30312 : mux21_ni port map ( Y=>nx30311, A0=>label_1_output_10, A1=>
      label_1_input_10, S0=>nx43401);
   ix17937 : mux21_ni port map ( Y=>nx17936, A0=>nx17932, A1=>
      label_1_input_state_machine_10, S0=>nx43057);
   ix30302 : mux21_ni port map ( Y=>nx30301, A0=>
      label_1_input_state_machine_10, A1=>data_in(10), S0=>nx43349);
   ix30272 : mux21_ni port map ( Y=>nx30271, A0=>label_1_output_8, A1=>
      label_1_input_8, S0=>nx43401);
   ix17873 : mux21_ni port map ( Y=>nx17872, A0=>nx17868, A1=>
      label_1_input_state_machine_8, S0=>nx43057);
   ix30262 : mux21_ni port map ( Y=>nx30261, A0=>
      label_1_input_state_machine_8, A1=>data_in(8), S0=>nx43349);
   ix30232 : mux21_ni port map ( Y=>nx30231, A0=>label_1_output_6, A1=>
      label_1_input_6, S0=>nx43401);
   ix17809 : mux21_ni port map ( Y=>nx17808, A0=>nx17804, A1=>
      label_1_input_state_machine_6, S0=>nx43057);
   ix30222 : mux21_ni port map ( Y=>nx30221, A0=>
      label_1_input_state_machine_6, A1=>data_in(6), S0=>nx43349);
   ix30192 : mux21_ni port map ( Y=>nx30191, A0=>label_1_output_4, A1=>
      label_1_input_4, S0=>nx43401);
   ix17745 : mux21_ni port map ( Y=>nx17744, A0=>nx17740, A1=>
      label_1_input_state_machine_4, S0=>nx43057);
   ix30182 : mux21_ni port map ( Y=>nx30181, A0=>
      label_1_input_state_machine_4, A1=>data_in(4), S0=>nx43351);
   ix30152 : mux21_ni port map ( Y=>nx30151, A0=>label_1_output_2, A1=>
      label_1_input_2, S0=>nx43403);
   ix17681 : mux21_ni port map ( Y=>nx17680, A0=>nx17676, A1=>
      label_1_input_state_machine_2, S0=>nx43057);
   ix30142 : mux21_ni port map ( Y=>nx30141, A0=>
      label_1_input_state_machine_2, A1=>data_in(2), S0=>nx43351);
   ix20822 : mux21_ni port map ( Y=>nx20821, A0=>label_1_output_0, A1=>
      label_1_input_0, S0=>nx43403);
   ix20812 : mux21_ni port map ( Y=>nx20811, A0=>
      label_1_input_state_machine_0, A1=>data_in(0), S0=>nx43351);
   ix20802 : mux21_ni port map ( Y=>nx20801, A0=>
      booth_booth_integration_output_0_12, A1=>nx2806, S0=>nx43123);
   ix2807 : mux21_ni port map ( Y=>nx2806, A0=>nx41807, A1=>
      booth_booth_integration_output_0_13, S0=>nx43131);
   ix20782 : mux21_ni port map ( Y=>nx20781, A0=>
      booth_booth_integration_output_0_13, A1=>nx2788, S0=>nx43123);
   ix2789 : mux21_ni port map ( Y=>nx2788, A0=>nx41803, A1=>
      booth_booth_integration_output_0_14, S0=>nx43131);
   ix20762 : mux21_ni port map ( Y=>nx20761, A0=>
      booth_booth_integration_output_0_14, A1=>nx2770, S0=>nx43123);
   ix2771 : mux21_ni port map ( Y=>nx2770, A0=>nx41799, A1=>
      booth_booth_integration_output_0_15, S0=>nx43131);
   ix20742 : mux21 port map ( Y=>nx20741, A0=>nx33280, A1=>nx32833, S0=>
      nx43123);
   ix20732 : mux21_ni port map ( Y=>nx20731, A0=>data_in(15), A1=>nx41795, 
      S0=>nx42983);
   ix1971 : or04 port map ( Y=>nx41733, A0=>nx36, A1=>nx32838, A2=>nx42273, 
      A3=>nx41381);
   ix32839 : or02 port map ( Y=>nx32838, A0=>rst, A1=>nx42257);
   ix20142 : mux21_ni port map ( Y=>nx20141, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_0, A1=>nx41721, S0=>nx42921
   );
   ix20128 : and02 port map ( Y=>nx20127, A0=>nx43463, A1=>
      booth_booth_integrtaion_0_shift_Reg_count_0);
   ix20322 : mux21_ni port map ( Y=>nx20321, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_9, A1=>nx41707, S0=>nx42921
   );
   ix20312 : mux21_ni port map ( Y=>nx20311, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_9, A1=>output_8_dup_12688, 
      S0=>nx43123);
   ix20302 : mux21_ni port map ( Y=>nx20301, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_8, A1=>output_8_dup_12688, 
      S0=>nx42921);
   ix20292 : mux21_ni port map ( Y=>nx20291, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_8, A1=>output_7_dup_12689, 
      S0=>nx43123);
   ix20282 : mux21_ni port map ( Y=>nx20281, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_7, A1=>output_7_dup_12689, 
      S0=>nx42921);
   ix20272 : mux21_ni port map ( Y=>nx20271, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_7, A1=>output_6_dup_12690, 
      S0=>nx43125);
   ix20262 : mux21_ni port map ( Y=>nx20261, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_6, A1=>output_6_dup_12690, 
      S0=>nx42921);
   ix20252 : mux21_ni port map ( Y=>nx20251, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_6, A1=>output_5_dup_12691, 
      S0=>nx43125);
   ix20242 : mux21_ni port map ( Y=>nx20241, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_5, A1=>output_5_dup_12691, 
      S0=>nx42921);
   ix20232 : mux21_ni port map ( Y=>nx20231, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_5, A1=>output_4_dup_12692, 
      S0=>nx43125);
   ix20222 : mux21_ni port map ( Y=>nx20221, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_4, A1=>output_4_dup_12692, 
      S0=>nx42923);
   ix20212 : mux21_ni port map ( Y=>nx20211, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_4, A1=>output_3_dup_12693, 
      S0=>nx43125);
   ix20202 : mux21_ni port map ( Y=>nx20201, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_3, A1=>output_3_dup_12693, 
      S0=>nx42923);
   ix20192 : mux21_ni port map ( Y=>nx20191, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_3, A1=>output_2_dup_12694, 
      S0=>nx43125);
   ix20182 : mux21_ni port map ( Y=>nx20181, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_2, A1=>output_2_dup_12694, 
      S0=>nx42923);
   ix20172 : mux21_ni port map ( Y=>nx20171, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_2, A1=>output_1_dup_12695, 
      S0=>nx43125);
   ix20162 : mux21_ni port map ( Y=>nx20161, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_1, A1=>output_1_dup_12695, 
      S0=>nx42923);
   ix20152 : mux21_ni port map ( Y=>nx20151, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_1, A1=>nx41721, S0=>nx43125
   );
   ix2199 : nand02 port map ( Y=>nx33023, A0=>nx32912, A1=>booth_output_0);
   ix32915 : or03 port map ( Y=>nx32914, A0=>nx32999, A1=>
      booth_booth_integrtaion_0_shift_reg_output_0, A2=>nx43463);
   ix20562 : mux21_ni port map ( Y=>nx20561, A0=>booth_output_0, A1=>nx2178, 
      S0=>nx43127);
   ix2179 : mux21_ni port map ( Y=>nx2178, A0=>nx41781, A1=>booth_output_1, 
      S0=>nx43133);
   ix20542 : mux21_ni port map ( Y=>nx20541, A0=>booth_output_1, A1=>nx2160, 
      S0=>nx43127);
   ix2161 : mux21_ni port map ( Y=>nx2160, A0=>nx41777, A1=>booth_output_2, 
      S0=>nx43133);
   ix20522 : mux21_ni port map ( Y=>nx20521, A0=>booth_output_2, A1=>nx2142, 
      S0=>nx43127);
   ix2143 : mux21_ni port map ( Y=>nx2142, A0=>nx41773, A1=>booth_output_3, 
      S0=>nx43133);
   ix20502 : mux21_ni port map ( Y=>nx20501, A0=>booth_output_3, A1=>nx2124, 
      S0=>nx43127);
   ix2125 : mux21_ni port map ( Y=>nx2124, A0=>nx41769, A1=>booth_output_4, 
      S0=>nx43133);
   ix20482 : mux21_ni port map ( Y=>nx20481, A0=>booth_output_4, A1=>nx2106, 
      S0=>nx43127);
   ix2107 : mux21_ni port map ( Y=>nx2106, A0=>nx41765, A1=>booth_output_5, 
      S0=>nx43133);
   ix20462 : mux21_ni port map ( Y=>nx20461, A0=>booth_output_5, A1=>nx2088, 
      S0=>nx43127);
   ix2089 : mux21_ni port map ( Y=>nx2088, A0=>nx41761, A1=>booth_output_6, 
      S0=>nx43133);
   ix20442 : mux21_ni port map ( Y=>nx20441, A0=>booth_output_6, A1=>nx2070, 
      S0=>nx43127);
   ix2071 : mux21_ni port map ( Y=>nx2070, A0=>nx41757, A1=>booth_output_7, 
      S0=>nx43133);
   ix20422 : mux21_ni port map ( Y=>nx20421, A0=>booth_output_7, A1=>nx2052, 
      S0=>nx43129);
   ix2053 : mux21_ni port map ( Y=>nx2052, A0=>nx41753, A1=>booth_output_8, 
      S0=>nx43135);
   ix20402 : mux21_ni port map ( Y=>nx20401, A0=>booth_output_8, A1=>nx2034, 
      S0=>nx43129);
   ix2035 : mux21_ni port map ( Y=>nx2034, A0=>nx41749, A1=>booth_output_9, 
      S0=>nx43135);
   ix20382 : mux21_ni port map ( Y=>nx20381, A0=>booth_output_9, A1=>nx2016, 
      S0=>nx43129);
   ix2017 : mux21_ni port map ( Y=>nx2016, A0=>nx41745, A1=>booth_output_10, 
      S0=>nx43135);
   ix20362 : mux21_ni port map ( Y=>nx20361, A0=>booth_output_10, A1=>nx1998, 
      S0=>nx43129);
   ix1999 : mux21_ni port map ( Y=>nx1998, A0=>nx41741, A1=>booth_output_11, 
      S0=>nx43135);
   ix20342 : mux21_ni port map ( Y=>nx20341, A0=>booth_output_11, A1=>nx1980, 
      S0=>nx43129);
   ix1981 : mux21_ni port map ( Y=>nx1980, A0=>nx41729, A1=>
      booth_booth_integration_output_0_12, S0=>nx43135);
   ix20332 : mux21_ni port map ( Y=>nx20331, A0=>data_in(11), A1=>nx41729, 
      S0=>nx42983);
   ix20352 : mux21_ni port map ( Y=>nx20351, A0=>data_in(10), A1=>nx41741, 
      S0=>nx42983);
   ix20372 : mux21_ni port map ( Y=>nx20371, A0=>data_in(9), A1=>nx41745, S0
      =>nx42983);
   ix20392 : mux21_ni port map ( Y=>nx20391, A0=>data_in(8), A1=>nx41749, S0
      =>nx42983);
   ix20412 : mux21_ni port map ( Y=>nx20411, A0=>data_in(7), A1=>nx41753, S0
      =>nx42983);
   ix20432 : mux21_ni port map ( Y=>nx20431, A0=>data_in(6), A1=>nx41757, S0
      =>nx42983);
   ix20452 : mux21_ni port map ( Y=>nx20451, A0=>data_in(5), A1=>nx41761, S0
      =>nx42985);
   ix20472 : mux21_ni port map ( Y=>nx20471, A0=>data_in(4), A1=>nx41765, S0
      =>nx42985);
   ix20492 : mux21_ni port map ( Y=>nx20491, A0=>data_in(3), A1=>nx41769, S0
      =>nx42985);
   ix20512 : mux21_ni port map ( Y=>nx20511, A0=>data_in(2), A1=>nx41773, S0
      =>nx42985);
   ix20532 : mux21_ni port map ( Y=>nx20531, A0=>data_in(1), A1=>nx41777, S0
      =>nx42985);
   ix20552 : mux21_ni port map ( Y=>nx20551, A0=>data_in(0), A1=>nx41781, S0
      =>nx42985);
   ix20722 : mux21_ni port map ( Y=>nx20721, A0=>
      booth_booth_integration_output_0_16, A1=>nx2728, S0=>nx43129);
   ix2729 : nor02ii port map ( Y=>nx2728, A0=>nx33005, A1=>nx43135);
   ix2205 : nor02ii port map ( Y=>nx2204, A0=>nx32907, A1=>
      booth_booth_integration_output_0_16);
   ix2723 : xor2 port map ( Y=>nx18195, A0=>nx33011, A1=>nx33273);
   ix33027 : or02 port map ( Y=>nx33026, A0=>nx32912, A1=>booth_output_0);
   ix2711 : xor2 port map ( Y=>nx18196, A0=>nx33031, A1=>nx42385);
   ix33045 : xor2 port map ( Y=>nx33044, A0=>nx33048, A1=>nx2276);
   ix33057 : nor02ii port map ( Y=>nx33056, A0=>nx2242, A1=>data_in(3));
   ix2687 : xor2 port map ( Y=>nx18198, A0=>nx33079, A1=>nx42387);
   ix20682 : mux21_ni port map ( Y=>nx20681, A0=>
      booth_booth_integration_output_0_20, A1=>nx2680, S0=>nx43129);
   ix2681 : nor02ii port map ( Y=>nx2680, A0=>nx33067, A1=>nx43135);
   ix2675 : xor2 port map ( Y=>nx18199, A0=>nx33084, A1=>nx33270);
   ix2663 : xor2 port map ( Y=>nx18200, A0=>nx33113, A1=>nx42389);
   ix20662 : mux21_ni port map ( Y=>nx20661, A0=>
      booth_booth_integration_output_0_22, A1=>nx2656, S0=>nx42379);
   ix2657 : nor02ii port map ( Y=>nx2656, A0=>nx33101, A1=>nx42383);
   ix2651 : xor2 port map ( Y=>nx18201, A0=>nx33118, A1=>nx33267);
   ix2639 : xor2 port map ( Y=>nx18203, A0=>nx33147, A1=>nx42391);
   ix20642 : mux21_ni port map ( Y=>nx20641, A0=>
      booth_booth_integration_output_0_24, A1=>nx2632, S0=>nx42379);
   ix2633 : nor02ii port map ( Y=>nx2632, A0=>nx33135, A1=>nx42383);
   ix2627 : xor2 port map ( Y=>nx18205, A0=>nx33152, A1=>nx33264);
   ix2615 : xor2 port map ( Y=>nx18207, A0=>nx33181, A1=>nx42393);
   ix20622 : mux21_ni port map ( Y=>nx20621, A0=>
      booth_booth_integration_output_0_26, A1=>nx2608, S0=>nx42379);
   ix2609 : nor02ii port map ( Y=>nx2608, A0=>nx33169, A1=>nx42383);
   ix2603 : xor2 port map ( Y=>nx18209, A0=>nx33186, A1=>nx33261);
   ix2591 : xor2 port map ( Y=>nx18210, A0=>nx33215, A1=>nx42395);
   ix20602 : mux21_ni port map ( Y=>nx20601, A0=>booth_output_28, A1=>nx2584, 
      S0=>nx42379);
   ix2585 : nor02ii port map ( Y=>nx2584, A0=>nx33203, A1=>nx42383);
   ix2579 : xor2 port map ( Y=>nx18211, A0=>nx33220, A1=>nx33258);
   ix2567 : xor2 port map ( Y=>nx18212, A0=>nx33236, A1=>nx42397);
   ix33252 : xor2 port map ( Y=>nx33251, A0=>nx33236, A1=>nx2552);
   ix2741 : nor02ii port map ( Y=>nx2740, A0=>nx2204, A1=>nx42383);
   ix20752 : mux21_ni port map ( Y=>nx20751, A0=>data_in(14), A1=>nx41799, 
      S0=>nx42985);
   ix20772 : mux21_ni port map ( Y=>nx20771, A0=>data_in(13), A1=>nx41803, 
      S0=>nx42987);
   ix20792 : mux21_ni port map ( Y=>nx20791, A0=>data_in(12), A1=>nx41807, 
      S0=>nx42987);
   ix33313 : nor02ii port map ( Y=>nx33312, A0=>sel_dst_0, A1=>nx43059);
   ix33316 : xnor2 port map ( Y=>nx33315, A0=>nx33289, A1=>nx33325);
   ix30132 : mux21_ni port map ( Y=>nx30131, A0=>label_1_output_1, A1=>
      label_1_input_1, S0=>nx43403);
   ix17649 : mux21_ni port map ( Y=>nx17648, A0=>nx17644, A1=>
      label_1_input_state_machine_1, S0=>nx43059);
   ix30122 : mux21_ni port map ( Y=>nx30121, A0=>
      label_1_input_state_machine_1, A1=>data_in(1), S0=>nx43351);
   ix33331 : xnor2 port map ( Y=>nx33330, A0=>nx33280, A1=>nx33340);
   ix30172 : mux21_ni port map ( Y=>nx30171, A0=>label_1_output_3, A1=>
      label_1_input_3, S0=>nx43403);
   ix17713 : mux21_ni port map ( Y=>nx17712, A0=>nx17708, A1=>
      label_1_input_state_machine_3, S0=>nx43059);
   ix30162 : mux21_ni port map ( Y=>nx30161, A0=>
      label_1_input_state_machine_3, A1=>data_in(3), S0=>nx43351);
   ix33342 : xor2 port map ( Y=>nx33341, A0=>nx33001, A1=>label_1_output_4);
   ix33346 : xnor2 port map ( Y=>nx33345, A0=>nx33011, A1=>nx33355);
   ix30212 : mux21_ni port map ( Y=>nx30211, A0=>label_1_output_5, A1=>
      label_1_input_5, S0=>nx43403);
   ix17777 : mux21_ni port map ( Y=>nx17776, A0=>nx17772, A1=>
      label_1_input_state_machine_5, S0=>nx43059);
   ix30202 : mux21_ni port map ( Y=>nx30201, A0=>
      label_1_input_state_machine_5, A1=>data_in(5), S0=>nx43351);
   ix33357 : xor2 port map ( Y=>nx33356, A0=>nx33031, A1=>label_1_output_6);
   ix33361 : xnor2 port map ( Y=>nx33360, A0=>nx33048, A1=>nx33370);
   ix30252 : mux21_ni port map ( Y=>nx30251, A0=>label_1_output_7, A1=>
      label_1_input_7, S0=>nx43403);
   ix17841 : mux21_ni port map ( Y=>nx17840, A0=>nx17836, A1=>
      label_1_input_state_machine_7, S0=>nx43059);
   ix30242 : mux21_ni port map ( Y=>nx30241, A0=>
      label_1_input_state_machine_7, A1=>data_in(7), S0=>nx43351);
   ix33372 : xor2 port map ( Y=>nx33371, A0=>nx33079, A1=>label_1_output_8);
   ix33376 : xnor2 port map ( Y=>nx33375, A0=>nx33084, A1=>nx33385);
   ix30292 : mux21_ni port map ( Y=>nx30291, A0=>label_1_output_9, A1=>
      label_1_input_9, S0=>nx43403);
   ix17905 : mux21_ni port map ( Y=>nx17904, A0=>nx17900, A1=>
      label_1_input_state_machine_9, S0=>nx43059);
   ix30282 : mux21_ni port map ( Y=>nx30281, A0=>
      label_1_input_state_machine_9, A1=>data_in(9), S0=>nx43353);
   ix33387 : xor2 port map ( Y=>nx33386, A0=>nx33113, A1=>label_1_output_10
   );
   ix33391 : xnor2 port map ( Y=>nx33390, A0=>nx33118, A1=>nx33400);
   ix30332 : mux21_ni port map ( Y=>nx30331, A0=>label_1_output_11, A1=>
      label_1_input_11, S0=>nx43405);
   ix17969 : mux21_ni port map ( Y=>nx17968, A0=>nx17964, A1=>
      label_1_input_state_machine_11, S0=>nx43059);
   ix30322 : mux21_ni port map ( Y=>nx30321, A0=>
      label_1_input_state_machine_11, A1=>data_in(11), S0=>nx43353);
   ix33402 : xor2 port map ( Y=>nx33401, A0=>nx33147, A1=>label_1_output_12
   );
   ix33406 : xnor2 port map ( Y=>nx33405, A0=>nx33152, A1=>nx33415);
   ix30372 : mux21_ni port map ( Y=>nx30371, A0=>label_1_output_13, A1=>
      label_1_input_13, S0=>nx43405);
   ix18033 : mux21_ni port map ( Y=>nx18032, A0=>nx18028, A1=>
      label_1_input_state_machine_13, S0=>nx42287);
   ix30362 : mux21_ni port map ( Y=>nx30361, A0=>
      label_1_input_state_machine_13, A1=>data_in(13), S0=>nx43353);
   ix33417 : xor2 port map ( Y=>nx33416, A0=>nx33181, A1=>label_1_output_14
   );
   ix20001 : xnor2 port map ( Y=>nx20000, A0=>nx33186, A1=>label_1_output_15
   );
   ix31592 : mux21_ni port map ( Y=>nx31591, A0=>nx18623, A1=>
      max_calc_ans1_15, S0=>nx42991);
   ix2867 : nand03 port map ( Y=>nx41821, A0=>nx43031, A1=>nx42925, A2=>
      nx42871);
   ix1783 : or02 port map ( Y=>nx1782, A0=>nx33436, A1=>nx43453);
   ix33445 : nor02ii port map ( Y=>nx33444, A0=>start_comp, A1=>nx31896);
   ix1733 : nor03_2x port map ( Y=>nx41575, A0=>nx33436, A1=>nx43137, A2=>
      nx42843);
   ix42842 : inv01 port map ( Y=>nx42843, A=>nx33447);
   ix33448 : and02 port map ( Y=>nx33447, A0=>max_calc_state_2, A1=>nx42925
   );
   ix33454 : xor2 port map ( Y=>nx33453, A0=>nx42217, A1=>nx34095);
   ix22822 : mux21_ni port map ( Y=>nx22821, A0=>label_10_output_15, A1=>
      label_10_input_15, S0=>nx43405);
   ix5917 : mux21_ni port map ( Y=>nx5916, A0=>nx5912, A1=>
      label_10_input_state_machine_15, S0=>nx43061);
   ix22812 : mux21_ni port map ( Y=>nx22811, A0=>
      label_10_input_state_machine_15, A1=>data_in(159), S0=>nx43353);
   ix22232 : mux21_ni port map ( Y=>nx22231, A0=>label_10_output_14, A1=>
      label_10_input_14, S0=>nx43405);
   ix5063 : mux21_ni port map ( Y=>nx5062, A0=>nx5058, A1=>
      label_10_input_state_machine_14, S0=>nx43061);
   ix21412 : mux21_ni port map ( Y=>nx21411, A0=>
      label_10_input_state_machine_14, A1=>data_in(158), S0=>nx43353);
   ix22202 : mux21_ni port map ( Y=>nx22201, A0=>label_10_output_12, A1=>
      label_10_input_12, S0=>nx43405);
   ix5005 : mux21_ni port map ( Y=>nx5004, A0=>nx5000, A1=>
      label_10_input_state_machine_12, S0=>nx43061);
   ix22192 : mux21_ni port map ( Y=>nx22191, A0=>
      label_10_input_state_machine_12, A1=>data_in(156), S0=>nx43353);
   ix22162 : mux21_ni port map ( Y=>nx22161, A0=>label_10_output_10, A1=>
      label_10_input_10, S0=>nx43405);
   ix4941 : mux21_ni port map ( Y=>nx4940, A0=>nx4936, A1=>
      label_10_input_state_machine_10, S0=>nx43061);
   ix22152 : mux21_ni port map ( Y=>nx22151, A0=>
      label_10_input_state_machine_10, A1=>data_in(154), S0=>nx43353);
   ix22122 : mux21_ni port map ( Y=>nx22121, A0=>label_10_output_8, A1=>
      label_10_input_8, S0=>nx43405);
   ix4877 : mux21_ni port map ( Y=>nx4876, A0=>nx4872, A1=>
      label_10_input_state_machine_8, S0=>nx43063);
   ix22112 : mux21_ni port map ( Y=>nx22111, A0=>
      label_10_input_state_machine_8, A1=>data_in(152), S0=>nx43355);
   ix22082 : mux21_ni port map ( Y=>nx22081, A0=>label_10_output_6, A1=>
      label_10_input_6, S0=>nx43407);
   ix4813 : mux21_ni port map ( Y=>nx4812, A0=>nx4808, A1=>
      label_10_input_state_machine_6, S0=>nx43063);
   ix22072 : mux21_ni port map ( Y=>nx22071, A0=>
      label_10_input_state_machine_6, A1=>data_in(150), S0=>nx43355);
   ix22042 : mux21_ni port map ( Y=>nx22041, A0=>label_10_output_4, A1=>
      label_10_input_4, S0=>nx43407);
   ix4749 : mux21_ni port map ( Y=>nx4748, A0=>nx4744, A1=>
      label_10_input_state_machine_4, S0=>nx43063);
   ix22032 : mux21_ni port map ( Y=>nx22031, A0=>
      label_10_input_state_machine_4, A1=>data_in(148), S0=>nx43355);
   ix22002 : mux21_ni port map ( Y=>nx22001, A0=>label_10_output_2, A1=>
      label_10_input_2, S0=>nx43407);
   ix4685 : mux21_ni port map ( Y=>nx4684, A0=>nx4680, A1=>
      label_10_input_state_machine_2, S0=>nx42287);
   ix21992 : mux21_ni port map ( Y=>nx21991, A0=>
      label_10_input_state_machine_2, A1=>data_in(146), S0=>nx43355);
   ix21962 : mux21_ni port map ( Y=>nx21961, A0=>label_10_output_0, A1=>
      label_10_input_0, S0=>nx43407);
   ix21952 : mux21_ni port map ( Y=>nx21951, A0=>
      label_10_input_state_machine_0, A1=>data_in(144), S0=>nx43355);
   ix21942 : mux21_ni port map ( Y=>nx21941, A0=>
      booth_booth_integration_output_9_12, A1=>nx4604, S0=>nx43163);
   ix4605 : mux21_ni port map ( Y=>nx4604, A0=>nx41807, A1=>
      booth_booth_integration_output_9_13, S0=>nx43171);
   ix21932 : mux21_ni port map ( Y=>nx21931, A0=>
      booth_booth_integration_output_9_13, A1=>nx4592, S0=>nx43163);
   ix4593 : mux21_ni port map ( Y=>nx4592, A0=>nx41803, A1=>
      booth_booth_integration_output_9_14, S0=>nx43171);
   ix21922 : mux21_ni port map ( Y=>nx21921, A0=>
      booth_booth_integration_output_9_14, A1=>nx4580, S0=>nx43163);
   ix4581 : mux21_ni port map ( Y=>nx4580, A0=>nx41799, A1=>
      booth_booth_integration_output_9_15, S0=>nx43171);
   ix21912 : mux21 port map ( Y=>nx21911, A0=>nx33982, A1=>nx33563, S0=>
      nx43163);
   ix21442 : mux21_ni port map ( Y=>nx21441, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_0, A1=>nx41879, S0=>nx42929
   );
   ix21428 : and02 port map ( Y=>nx21427, A0=>nx43471, A1=>
      booth_booth_integrtaion_9_shift_Reg_count_0);
   ix21622 : mux21_ni port map ( Y=>nx21621, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_9, A1=>nx41865, S0=>nx42929
   );
   ix21612 : mux21_ni port map ( Y=>nx21611, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_9, A1=>output_8_dup_12940, 
      S0=>nx43163);
   ix21602 : mux21_ni port map ( Y=>nx21601, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_8, A1=>output_8_dup_12940, 
      S0=>nx42929);
   ix21592 : mux21_ni port map ( Y=>nx21591, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_8, A1=>output_7_dup_12941, 
      S0=>nx43163);
   ix21582 : mux21_ni port map ( Y=>nx21581, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_7, A1=>output_7_dup_12941, 
      S0=>nx42929);
   ix21572 : mux21_ni port map ( Y=>nx21571, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_7, A1=>output_6_dup_12942, 
      S0=>nx43165);
   ix21562 : mux21_ni port map ( Y=>nx21561, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_6, A1=>output_6_dup_12942, 
      S0=>nx42929);
   ix21552 : mux21_ni port map ( Y=>nx21551, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_6, A1=>output_5_dup_12943, 
      S0=>nx43165);
   ix21542 : mux21_ni port map ( Y=>nx21541, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_5, A1=>output_5_dup_12943, 
      S0=>nx42929);
   ix21532 : mux21_ni port map ( Y=>nx21531, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_5, A1=>output_4_dup_12944, 
      S0=>nx43165);
   ix21522 : mux21_ni port map ( Y=>nx21521, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_4, A1=>output_4_dup_12944, 
      S0=>nx42931);
   ix21512 : mux21_ni port map ( Y=>nx21511, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_4, A1=>output_3_dup_12945, 
      S0=>nx43165);
   ix21502 : mux21_ni port map ( Y=>nx21501, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_3, A1=>output_3_dup_12945, 
      S0=>nx42931);
   ix21492 : mux21_ni port map ( Y=>nx21491, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_3, A1=>output_2_dup_12946, 
      S0=>nx43165);
   ix21482 : mux21_ni port map ( Y=>nx21481, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_2, A1=>output_2_dup_12946, 
      S0=>nx42931);
   ix21472 : mux21_ni port map ( Y=>nx21471, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_2, A1=>output_1_dup_12947, 
      S0=>nx43165);
   ix21462 : mux21_ni port map ( Y=>nx21461, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_1, A1=>output_1_dup_12947, 
      S0=>nx42931);
   ix21452 : mux21_ni port map ( Y=>nx21451, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_1, A1=>nx41879, S0=>nx43165
   );
   ix4021 : nand02 port map ( Y=>nx33709, A0=>nx33636, A1=>
      booth_output_0_dup_12282);
   ix33639 : or03 port map ( Y=>nx33638, A0=>nx33687, A1=>
      booth_booth_integrtaion_9_shift_reg_output_0, A2=>nx43471);
   ix21742 : mux21_ni port map ( Y=>nx21741, A0=>booth_output_0_dup_12282, 
      A1=>nx4000, S0=>nx43167);
   ix4001 : mux21_ni port map ( Y=>nx4000, A0=>nx41781, A1=>
      booth_output_1_dup_12281, S0=>nx43173);
   ix21732 : mux21_ni port map ( Y=>nx21731, A0=>booth_output_1_dup_12281, 
      A1=>nx3988, S0=>nx43167);
   ix3989 : mux21_ni port map ( Y=>nx3988, A0=>nx41777, A1=>
      booth_output_2_dup_12280, S0=>nx43173);
   ix21722 : mux21_ni port map ( Y=>nx21721, A0=>booth_output_2_dup_12280, 
      A1=>nx3976, S0=>nx43167);
   ix3977 : mux21_ni port map ( Y=>nx3976, A0=>nx41773, A1=>
      booth_output_3_dup_12279, S0=>nx43173);
   ix21712 : mux21_ni port map ( Y=>nx21711, A0=>booth_output_3_dup_12279, 
      A1=>nx3964, S0=>nx43167);
   ix3965 : mux21_ni port map ( Y=>nx3964, A0=>nx41769, A1=>
      booth_output_4_dup_12278, S0=>nx43173);
   ix21702 : mux21_ni port map ( Y=>nx21701, A0=>booth_output_4_dup_12278, 
      A1=>nx3952, S0=>nx43167);
   ix3953 : mux21_ni port map ( Y=>nx3952, A0=>nx41765, A1=>
      booth_output_5_dup_12277, S0=>nx43173);
   ix21692 : mux21_ni port map ( Y=>nx21691, A0=>booth_output_5_dup_12277, 
      A1=>nx3940, S0=>nx43167);
   ix3941 : mux21_ni port map ( Y=>nx3940, A0=>nx41761, A1=>
      booth_output_6_dup_12276, S0=>nx43173);
   ix21682 : mux21_ni port map ( Y=>nx21681, A0=>booth_output_6_dup_12276, 
      A1=>nx3928, S0=>nx43167);
   ix3929 : mux21_ni port map ( Y=>nx3928, A0=>nx41757, A1=>
      booth_output_7_dup_12275, S0=>nx43173);
   ix21672 : mux21_ni port map ( Y=>nx21671, A0=>booth_output_7_dup_12275, 
      A1=>nx3916, S0=>nx43169);
   ix3917 : mux21_ni port map ( Y=>nx3916, A0=>nx41753, A1=>
      booth_output_8_dup_12274, S0=>nx43175);
   ix21662 : mux21_ni port map ( Y=>nx21661, A0=>booth_output_8_dup_12274, 
      A1=>nx3904, S0=>nx43169);
   ix3905 : mux21_ni port map ( Y=>nx3904, A0=>nx41749, A1=>
      booth_output_9_dup_12273, S0=>nx43175);
   ix21652 : mux21_ni port map ( Y=>nx21651, A0=>booth_output_9_dup_12273, 
      A1=>nx3892, S0=>nx43169);
   ix3893 : mux21_ni port map ( Y=>nx3892, A0=>nx41745, A1=>
      booth_output_10_dup_12272, S0=>nx43175);
   ix21642 : mux21_ni port map ( Y=>nx21641, A0=>booth_output_10_dup_12272, 
      A1=>nx3880, S0=>nx43169);
   ix3881 : mux21_ni port map ( Y=>nx3880, A0=>nx41741, A1=>
      booth_output_11_dup_12271, S0=>nx43175);
   ix21632 : mux21_ni port map ( Y=>nx21631, A0=>booth_output_11_dup_12271, 
      A1=>nx3868, S0=>nx43169);
   ix3869 : mux21_ni port map ( Y=>nx3868, A0=>nx41729, A1=>
      booth_booth_integration_output_9_12, S0=>nx43175);
   ix21902 : mux21_ni port map ( Y=>nx21901, A0=>
      booth_booth_integration_output_9_16, A1=>nx4550, S0=>nx43169);
   ix4551 : nor02ii port map ( Y=>nx4550, A0=>nx33693, A1=>nx43175);
   ix4027 : nor02ii port map ( Y=>nx4026, A0=>nx33631, A1=>
      booth_booth_integration_output_9_16);
   ix4545 : xor2 port map ( Y=>nx18239, A0=>nx33699, A1=>nx33975);
   ix33715 : or02 port map ( Y=>nx33714, A0=>nx33636, A1=>
      booth_output_0_dup_12282);
   ix4533 : xor2 port map ( Y=>nx18241, A0=>nx33719, A1=>nx42471);
   ix33735 : xor2 port map ( Y=>nx33734, A0=>nx33738, A1=>nx4098);
   ix33747 : nor02ii port map ( Y=>nx33746, A0=>nx4064, A1=>data_in(147));
   ix4509 : xor2 port map ( Y=>nx18243, A0=>nx33771, A1=>nx42473);
   ix21862 : mux21_ni port map ( Y=>nx21861, A0=>
      booth_booth_integration_output_9_20, A1=>nx4502, S0=>nx43169);
   ix4503 : nor02ii port map ( Y=>nx4502, A0=>nx33757, A1=>nx43175);
   ix4497 : xor2 port map ( Y=>nx18244, A0=>nx33776, A1=>nx33972);
   ix4485 : xor2 port map ( Y=>nx18245, A0=>nx33807, A1=>nx42475);
   ix21842 : mux21_ni port map ( Y=>nx21841, A0=>
      booth_booth_integration_output_9_22, A1=>nx4478, S0=>nx42465);
   ix4479 : nor02ii port map ( Y=>nx4478, A0=>nx33793, A1=>nx42469);
   ix4473 : xor2 port map ( Y=>nx18246, A0=>nx33812, A1=>nx33969);
   ix4461 : xor2 port map ( Y=>nx18247, A0=>nx33843, A1=>nx42477);
   ix21822 : mux21_ni port map ( Y=>nx21821, A0=>
      booth_booth_integration_output_9_24, A1=>nx4454, S0=>nx42465);
   ix4455 : nor02ii port map ( Y=>nx4454, A0=>nx33829, A1=>nx42469);
   ix4449 : xor2 port map ( Y=>nx18249, A0=>nx33848, A1=>nx33966);
   ix4437 : xor2 port map ( Y=>nx18251, A0=>nx33879, A1=>nx42479);
   ix21802 : mux21_ni port map ( Y=>nx21801, A0=>
      booth_booth_integration_output_9_26, A1=>nx4430, S0=>nx42465);
   ix4431 : nor02ii port map ( Y=>nx4430, A0=>nx33865, A1=>nx42469);
   ix4425 : xor2 port map ( Y=>nx18253, A0=>nx33884, A1=>nx33963);
   ix4413 : xor2 port map ( Y=>nx18254, A0=>nx33915, A1=>nx42481);
   ix21782 : mux21_ni port map ( Y=>nx21781, A0=>booth_output_28_dup_12270, 
      A1=>nx4406, S0=>nx42465);
   ix4407 : nor02ii port map ( Y=>nx4406, A0=>nx33901, A1=>nx42469);
   ix4401 : xor2 port map ( Y=>nx18255, A0=>nx33920, A1=>nx33960);
   ix4389 : xor2 port map ( Y=>nx18256, A0=>nx33936, A1=>nx42483);
   ix33954 : xor2 port map ( Y=>nx33953, A0=>nx33936, A1=>nx4374);
   ix4563 : nor02ii port map ( Y=>nx4562, A0=>nx4026, A1=>nx42469);
   ix33990 : xnor2 port map ( Y=>nx33989, A0=>nx33985, A1=>nx33999);
   ix21982 : mux21_ni port map ( Y=>nx21981, A0=>label_10_output_1, A1=>
      label_10_input_1, S0=>nx43407);
   ix4653 : mux21_ni port map ( Y=>nx4652, A0=>nx4648, A1=>
      label_10_input_state_machine_1, S0=>nx42287);
   ix21972 : mux21_ni port map ( Y=>nx21971, A0=>
      label_10_input_state_machine_1, A1=>data_in(145), S0=>nx43355);
   ix34005 : xnor2 port map ( Y=>nx34004, A0=>nx33982, A1=>nx34014);
   ix22022 : mux21_ni port map ( Y=>nx22021, A0=>label_10_output_3, A1=>
      label_10_input_3, S0=>nx43407);
   ix4717 : mux21_ni port map ( Y=>nx4716, A0=>nx4712, A1=>
      label_10_input_state_machine_3, S0=>nx43063);
   ix22012 : mux21_ni port map ( Y=>nx22011, A0=>
      label_10_input_state_machine_3, A1=>data_in(147), S0=>nx43355);
   ix34016 : xor2 port map ( Y=>nx34015, A0=>nx33689, A1=>label_10_output_4
   );
   ix34020 : xnor2 port map ( Y=>nx34019, A0=>nx33699, A1=>nx34029);
   ix22062 : mux21_ni port map ( Y=>nx22061, A0=>label_10_output_5, A1=>
      label_10_input_5, S0=>nx43407);
   ix4781 : mux21_ni port map ( Y=>nx4780, A0=>nx4776, A1=>
      label_10_input_state_machine_5, S0=>nx43063);
   ix22052 : mux21_ni port map ( Y=>nx22051, A0=>
      label_10_input_state_machine_5, A1=>data_in(149), S0=>nx43357);
   ix34031 : xor2 port map ( Y=>nx34030, A0=>nx33719, A1=>label_10_output_6
   );
   ix34035 : xnor2 port map ( Y=>nx34034, A0=>nx33738, A1=>nx34044);
   ix22102 : mux21_ni port map ( Y=>nx22101, A0=>label_10_output_7, A1=>
      label_10_input_7, S0=>nx43409);
   ix4845 : mux21_ni port map ( Y=>nx4844, A0=>nx4840, A1=>
      label_10_input_state_machine_7, S0=>nx43063);
   ix22092 : mux21_ni port map ( Y=>nx22091, A0=>
      label_10_input_state_machine_7, A1=>data_in(151), S0=>nx43357);
   ix34046 : xor2 port map ( Y=>nx34045, A0=>nx33771, A1=>label_10_output_8
   );
   ix34050 : xnor2 port map ( Y=>nx34049, A0=>nx33776, A1=>nx34059);
   ix22142 : mux21_ni port map ( Y=>nx22141, A0=>label_10_output_9, A1=>
      label_10_input_9, S0=>nx43409);
   ix4909 : mux21_ni port map ( Y=>nx4908, A0=>nx4904, A1=>
      label_10_input_state_machine_9, S0=>nx43063);
   ix22132 : mux21_ni port map ( Y=>nx22131, A0=>
      label_10_input_state_machine_9, A1=>data_in(153), S0=>nx43357);
   ix34061 : xor2 port map ( Y=>nx34060, A0=>nx33807, A1=>label_10_output_10
   );
   ix34065 : xnor2 port map ( Y=>nx34064, A0=>nx33812, A1=>nx34074);
   ix22182 : mux21_ni port map ( Y=>nx22181, A0=>label_10_output_11, A1=>
      label_10_input_11, S0=>nx43409);
   ix4973 : mux21_ni port map ( Y=>nx4972, A0=>nx4968, A1=>
      label_10_input_state_machine_11, S0=>nx43065);
   ix22172 : mux21_ni port map ( Y=>nx22171, A0=>
      label_10_input_state_machine_11, A1=>data_in(155), S0=>nx43357);
   ix34076 : xor2 port map ( Y=>nx34075, A0=>nx33843, A1=>label_10_output_12
   );
   ix34080 : xnor2 port map ( Y=>nx34079, A0=>nx33848, A1=>nx34089);
   ix22222 : mux21_ni port map ( Y=>nx22221, A0=>label_10_output_13, A1=>
      label_10_input_13, S0=>nx43409);
   ix5037 : mux21_ni port map ( Y=>nx5036, A0=>nx5032, A1=>
      label_10_input_state_machine_13, S0=>nx43065);
   ix22212 : mux21_ni port map ( Y=>nx22211, A0=>
      label_10_input_state_machine_13, A1=>data_in(157), S0=>nx43357);
   ix34091 : xor2 port map ( Y=>nx34090, A0=>nx33879, A1=>label_10_output_14
   );
   ix5911 : xnor2 port map ( Y=>nx5910, A0=>nx33884, A1=>label_10_output_15
   );
   ix31802 : mux21_ni port map ( Y=>nx31801, A0=>nx42213, A1=>nx18603, S0=>
      nx43335);
   ix18133 : mux21_ni port map ( Y=>nx18603, A0=>
      max_calc_comparator_first_inp2_14, A1=>
      max_calc_comparator_first_inp1_14, S0=>nx43025);
   ix30422 : mux21_ni port map ( Y=>nx30421, A0=>
      max_calc_comparator_first_inp1_14, A1=>nx18118, S0=>nx43391);
   ix18119 : mux21_ni port map ( Y=>nx18118, A0=>nx18114, A1=>nx18082, S0=>
      nx43031);
   ix18083 : mux21_ni port map ( Y=>nx18082, A0=>max_calc_ans1_14, A1=>
      label_1_output_14, S0=>nx43137);
   ix30392 : mux21_ni port map ( Y=>nx30391, A0=>nx18603, A1=>
      max_calc_ans1_14, S0=>nx42991);
   ix18115 : mux21_ni port map ( Y=>nx18114, A0=>max_calc_ans5_14, A1=>
      max_calc_ans6_14, S0=>nx43137);
   ix30402 : mux21_ni port map ( Y=>nx30401, A0=>max_calc_ans6_14, A1=>
      nx18603, S0=>nx43179);
   ix34113 : nor02ii port map ( Y=>nx42485, A0=>nx43203, A1=>nx34114);
   ix34115 : and02 port map ( Y=>nx34114, A0=>nx33436, A1=>nx43137);
   ix30412 : mux21_ni port map ( Y=>nx30411, A0=>max_calc_ans5_14, A1=>
      nx18104, S0=>nx42871);
   ix18105 : mux21 port map ( Y=>nx18104, A0=>nx34760, A1=>nx34125, S0=>
      nx43001);
   ix22522 : mux21_ni port map ( Y=>nx22521, A0=>label_9_output_14, A1=>
      label_9_input_14, S0=>nx43409);
   ix5513 : mux21_ni port map ( Y=>nx5512, A0=>nx5508, A1=>
      label_9_input_state_machine_14, S0=>nx43065);
   ix22252 : mux21_ni port map ( Y=>nx22251, A0=>
      label_9_input_state_machine_14, A1=>data_in(142), S0=>nx43357);
   ix22492 : mux21_ni port map ( Y=>nx22491, A0=>label_9_output_12, A1=>
      label_9_input_12, S0=>nx43409);
   ix5455 : mux21_ni port map ( Y=>nx5454, A0=>nx5450, A1=>
      label_9_input_state_machine_12, S0=>nx43065);
   ix22482 : mux21_ni port map ( Y=>nx22481, A0=>
      label_9_input_state_machine_12, A1=>data_in(140), S0=>nx43357);
   ix22452 : mux21_ni port map ( Y=>nx22451, A0=>label_9_output_10, A1=>
      label_9_input_10, S0=>nx43409);
   ix5391 : mux21_ni port map ( Y=>nx5390, A0=>nx5386, A1=>
      label_9_input_state_machine_10, S0=>nx43065);
   ix22442 : mux21_ni port map ( Y=>nx22441, A0=>
      label_9_input_state_machine_10, A1=>data_in(138), S0=>nx43359);
   ix22412 : mux21_ni port map ( Y=>nx22411, A0=>label_9_output_8, A1=>
      label_9_input_8, S0=>nx43411);
   ix5327 : mux21_ni port map ( Y=>nx5326, A0=>nx5322, A1=>
      label_9_input_state_machine_8, S0=>nx43065);
   ix22402 : mux21_ni port map ( Y=>nx22401, A0=>
      label_9_input_state_machine_8, A1=>data_in(136), S0=>nx43359);
   ix22372 : mux21_ni port map ( Y=>nx22371, A0=>label_9_output_6, A1=>
      label_9_input_6, S0=>nx43411);
   ix5263 : mux21_ni port map ( Y=>nx5262, A0=>nx5258, A1=>
      label_9_input_state_machine_6, S0=>nx43065);
   ix22362 : mux21_ni port map ( Y=>nx22361, A0=>
      label_9_input_state_machine_6, A1=>data_in(134), S0=>nx43359);
   ix22332 : mux21_ni port map ( Y=>nx22331, A0=>label_9_output_4, A1=>
      label_9_input_4, S0=>nx43411);
   ix5199 : mux21_ni port map ( Y=>nx5198, A0=>nx5194, A1=>
      label_9_input_state_machine_4, S0=>nx43067);
   ix22322 : mux21_ni port map ( Y=>nx22321, A0=>
      label_9_input_state_machine_4, A1=>data_in(132), S0=>nx43359);
   ix22292 : mux21_ni port map ( Y=>nx22291, A0=>label_9_output_2, A1=>
      label_9_input_2, S0=>nx43411);
   ix5135 : mux21_ni port map ( Y=>nx5134, A0=>nx5130, A1=>
      label_9_input_state_machine_2, S0=>nx43067);
   ix22282 : mux21_ni port map ( Y=>nx22281, A0=>
      label_9_input_state_machine_2, A1=>data_in(130), S0=>nx43359);
   ix21392 : mux21_ni port map ( Y=>nx21391, A0=>label_9_output_0, A1=>
      label_9_input_0, S0=>nx43411);
   ix21382 : mux21_ni port map ( Y=>nx21381, A0=>
      label_9_input_state_machine_0, A1=>data_in(128), S0=>nx43359);
   ix21372 : mux21_ni port map ( Y=>nx21371, A0=>
      booth_booth_integration_output_8_12, A1=>nx3724, S0=>nx43189);
   ix3725 : mux21_ni port map ( Y=>nx3724, A0=>nx41807, A1=>
      booth_booth_integration_output_8_13, S0=>nx43197);
   ix21362 : mux21_ni port map ( Y=>nx21361, A0=>
      booth_booth_integration_output_8_13, A1=>nx3712, S0=>nx43189);
   ix3713 : mux21_ni port map ( Y=>nx3712, A0=>nx41803, A1=>
      booth_booth_integration_output_8_14, S0=>nx43197);
   ix21352 : mux21_ni port map ( Y=>nx21351, A0=>
      booth_booth_integration_output_8_14, A1=>nx3700, S0=>nx43189);
   ix3701 : mux21_ni port map ( Y=>nx3700, A0=>nx41799, A1=>
      booth_booth_integration_output_8_15, S0=>nx43197);
   ix21342 : mux21 port map ( Y=>nx21341, A0=>nx34647, A1=>nx34228, S0=>
      nx43189);
   ix20872 : mux21_ni port map ( Y=>nx20871, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_0, A1=>nx41847, S0=>nx42933
   );
   ix20858 : and02 port map ( Y=>nx20857, A0=>nx43467, A1=>
      booth_booth_integrtaion_8_shift_Reg_count_0);
   ix21052 : mux21_ni port map ( Y=>nx21051, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_9, A1=>nx41833, S0=>nx42933
   );
   ix21042 : mux21_ni port map ( Y=>nx21041, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_9, A1=>output_8_dup_12912, 
      S0=>nx43189);
   ix21032 : mux21_ni port map ( Y=>nx21031, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_8, A1=>output_8_dup_12912, 
      S0=>nx42933);
   ix21022 : mux21_ni port map ( Y=>nx21021, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_8, A1=>output_7_dup_12913, 
      S0=>nx43189);
   ix21012 : mux21_ni port map ( Y=>nx21011, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_7, A1=>output_7_dup_12913, 
      S0=>nx42933);
   ix21002 : mux21_ni port map ( Y=>nx21001, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_7, A1=>output_6_dup_12914, 
      S0=>nx43191);
   ix20992 : mux21_ni port map ( Y=>nx20991, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_6, A1=>output_6_dup_12914, 
      S0=>nx42933);
   ix20982 : mux21_ni port map ( Y=>nx20981, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_6, A1=>output_5_dup_12915, 
      S0=>nx43191);
   ix20972 : mux21_ni port map ( Y=>nx20971, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_5, A1=>output_5_dup_12915, 
      S0=>nx42933);
   ix20962 : mux21_ni port map ( Y=>nx20961, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_5, A1=>output_4_dup_12916, 
      S0=>nx43191);
   ix20952 : mux21_ni port map ( Y=>nx20951, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_4, A1=>output_4_dup_12916, 
      S0=>nx42935);
   ix20942 : mux21_ni port map ( Y=>nx20941, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_4, A1=>output_3_dup_12917, 
      S0=>nx43191);
   ix20932 : mux21_ni port map ( Y=>nx20931, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_3, A1=>output_3_dup_12917, 
      S0=>nx42935);
   ix20922 : mux21_ni port map ( Y=>nx20921, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_3, A1=>output_2_dup_12918, 
      S0=>nx43191);
   ix20912 : mux21_ni port map ( Y=>nx20911, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_2, A1=>output_2_dup_12918, 
      S0=>nx42935);
   ix20902 : mux21_ni port map ( Y=>nx20901, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_2, A1=>output_1_dup_12919, 
      S0=>nx43191);
   ix20892 : mux21_ni port map ( Y=>nx20891, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_1, A1=>output_1_dup_12919, 
      S0=>nx42935);
   ix20882 : mux21_ni port map ( Y=>nx20881, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_1, A1=>nx41847, S0=>nx43191
   );
   ix3141 : nand02 port map ( Y=>nx34374, A0=>nx34301, A1=>
      booth_output_0_dup_12263);
   ix34304 : or03 port map ( Y=>nx34303, A0=>nx34352, A1=>
      booth_booth_integrtaion_8_shift_reg_output_0, A2=>nx43467);
   ix21172 : mux21_ni port map ( Y=>nx21171, A0=>booth_output_0_dup_12263, 
      A1=>nx3120, S0=>nx43193);
   ix3121 : mux21_ni port map ( Y=>nx3120, A0=>nx41781, A1=>
      booth_output_1_dup_12262, S0=>nx43199);
   ix21162 : mux21_ni port map ( Y=>nx21161, A0=>booth_output_1_dup_12262, 
      A1=>nx3108, S0=>nx43193);
   ix3109 : mux21_ni port map ( Y=>nx3108, A0=>nx41777, A1=>
      booth_output_2_dup_12261, S0=>nx43199);
   ix21152 : mux21_ni port map ( Y=>nx21151, A0=>booth_output_2_dup_12261, 
      A1=>nx3096, S0=>nx43193);
   ix3097 : mux21_ni port map ( Y=>nx3096, A0=>nx41773, A1=>
      booth_output_3_dup_12260, S0=>nx43199);
   ix21142 : mux21_ni port map ( Y=>nx21141, A0=>booth_output_3_dup_12260, 
      A1=>nx3084, S0=>nx43193);
   ix3085 : mux21_ni port map ( Y=>nx3084, A0=>nx41769, A1=>
      booth_output_4_dup_12259, S0=>nx43199);
   ix21132 : mux21_ni port map ( Y=>nx21131, A0=>booth_output_4_dup_12259, 
      A1=>nx3072, S0=>nx43193);
   ix3073 : mux21_ni port map ( Y=>nx3072, A0=>nx41765, A1=>
      booth_output_5_dup_12258, S0=>nx43199);
   ix21122 : mux21_ni port map ( Y=>nx21121, A0=>booth_output_5_dup_12258, 
      A1=>nx3060, S0=>nx43193);
   ix3061 : mux21_ni port map ( Y=>nx3060, A0=>nx41761, A1=>
      booth_output_6_dup_12257, S0=>nx43199);
   ix21112 : mux21_ni port map ( Y=>nx21111, A0=>booth_output_6_dup_12257, 
      A1=>nx3048, S0=>nx43193);
   ix3049 : mux21_ni port map ( Y=>nx3048, A0=>nx41757, A1=>
      booth_output_7_dup_12256, S0=>nx43199);
   ix21102 : mux21_ni port map ( Y=>nx21101, A0=>booth_output_7_dup_12256, 
      A1=>nx3036, S0=>nx43195);
   ix3037 : mux21_ni port map ( Y=>nx3036, A0=>nx41753, A1=>
      booth_output_8_dup_12255, S0=>nx43201);
   ix21092 : mux21_ni port map ( Y=>nx21091, A0=>booth_output_8_dup_12255, 
      A1=>nx3024, S0=>nx43195);
   ix3025 : mux21_ni port map ( Y=>nx3024, A0=>nx41749, A1=>
      booth_output_9_dup_12254, S0=>nx43201);
   ix21082 : mux21_ni port map ( Y=>nx21081, A0=>booth_output_9_dup_12254, 
      A1=>nx3012, S0=>nx43195);
   ix3013 : mux21_ni port map ( Y=>nx3012, A0=>nx41745, A1=>
      booth_output_10_dup_12253, S0=>nx43201);
   ix21072 : mux21_ni port map ( Y=>nx21071, A0=>booth_output_10_dup_12253, 
      A1=>nx3000, S0=>nx43195);
   ix3001 : mux21_ni port map ( Y=>nx3000, A0=>nx41741, A1=>
      booth_output_11_dup_12252, S0=>nx43201);
   ix21062 : mux21_ni port map ( Y=>nx21061, A0=>booth_output_11_dup_12252, 
      A1=>nx2988, S0=>nx43195);
   ix2989 : mux21_ni port map ( Y=>nx2988, A0=>nx41729, A1=>
      booth_booth_integration_output_8_12, S0=>nx43201);
   ix21332 : mux21_ni port map ( Y=>nx21331, A0=>
      booth_booth_integration_output_8_16, A1=>nx3670, S0=>nx43195);
   ix3671 : nor02ii port map ( Y=>nx3670, A0=>nx34358, A1=>nx43201);
   ix3147 : nor02ii port map ( Y=>nx3146, A0=>nx34296, A1=>
      booth_booth_integration_output_8_16);
   ix3665 : xor2 port map ( Y=>nx18215, A0=>nx34364, A1=>nx34640);
   ix34380 : or02 port map ( Y=>nx34379, A0=>nx34301, A1=>
      booth_output_0_dup_12263);
   ix3653 : xor2 port map ( Y=>nx18217, A0=>nx34384, A1=>nx42509);
   ix34400 : xor2 port map ( Y=>nx34399, A0=>nx34403, A1=>nx3218);
   ix34412 : nor02ii port map ( Y=>nx34411, A0=>nx3184, A1=>data_in(131));
   ix3629 : xor2 port map ( Y=>nx18221, A0=>nx34436, A1=>nx42511);
   ix21292 : mux21_ni port map ( Y=>nx21291, A0=>
      booth_booth_integration_output_8_20, A1=>nx3622, S0=>nx43195);
   ix3623 : nor02ii port map ( Y=>nx3622, A0=>nx34422, A1=>nx43201);
   ix3617 : xor2 port map ( Y=>nx18223, A0=>nx34441, A1=>nx34637);
   ix3605 : xor2 port map ( Y=>nx18225, A0=>nx34472, A1=>nx42513);
   ix21272 : mux21_ni port map ( Y=>nx21271, A0=>
      booth_booth_integration_output_8_22, A1=>nx3598, S0=>nx42503);
   ix3599 : nor02ii port map ( Y=>nx3598, A0=>nx34458, A1=>nx42507);
   ix3593 : xor2 port map ( Y=>nx18227, A0=>nx34477, A1=>nx34634);
   ix3581 : xor2 port map ( Y=>nx18228, A0=>nx34508, A1=>nx42515);
   ix21252 : mux21_ni port map ( Y=>nx21251, A0=>
      booth_booth_integration_output_8_24, A1=>nx3574, S0=>nx42503);
   ix3575 : nor02ii port map ( Y=>nx3574, A0=>nx34494, A1=>nx42507);
   ix3569 : xor2 port map ( Y=>nx18229, A0=>nx34513, A1=>nx34631);
   ix3557 : xor2 port map ( Y=>nx18230, A0=>nx34544, A1=>nx42517);
   ix21232 : mux21_ni port map ( Y=>nx21231, A0=>
      booth_booth_integration_output_8_26, A1=>nx3550, S0=>nx42503);
   ix3551 : nor02ii port map ( Y=>nx3550, A0=>nx34530, A1=>nx42507);
   ix3545 : xor2 port map ( Y=>nx18231, A0=>nx34549, A1=>nx34628);
   ix3533 : xor2 port map ( Y=>nx18232, A0=>nx34580, A1=>nx42519);
   ix21212 : mux21_ni port map ( Y=>nx21211, A0=>booth_output_28_dup_12251, 
      A1=>nx3526, S0=>nx42503);
   ix3527 : nor02ii port map ( Y=>nx3526, A0=>nx34566, A1=>nx42507);
   ix3521 : xor2 port map ( Y=>nx18233, A0=>nx34585, A1=>nx34625);
   ix3509 : xor2 port map ( Y=>nx18235, A0=>nx34601, A1=>nx42521);
   ix34619 : xor2 port map ( Y=>nx34618, A0=>nx34601, A1=>nx3494);
   ix3683 : nor02ii port map ( Y=>nx3682, A0=>nx3146, A1=>nx42507);
   ix34655 : xnor2 port map ( Y=>nx34654, A0=>nx34650, A1=>nx34664);
   ix22272 : mux21_ni port map ( Y=>nx22271, A0=>label_9_output_1, A1=>
      label_9_input_1, S0=>nx43411);
   ix5103 : mux21_ni port map ( Y=>nx5102, A0=>nx5098, A1=>
      label_9_input_state_machine_1, S0=>nx43067);
   ix22262 : mux21_ni port map ( Y=>nx22261, A0=>
      label_9_input_state_machine_1, A1=>data_in(129), S0=>nx43359);
   ix34670 : xnor2 port map ( Y=>nx34669, A0=>nx34647, A1=>nx34679);
   ix22312 : mux21_ni port map ( Y=>nx22311, A0=>label_9_output_3, A1=>
      label_9_input_3, S0=>nx43411);
   ix5167 : mux21_ni port map ( Y=>nx5166, A0=>nx5162, A1=>
      label_9_input_state_machine_3, S0=>nx43067);
   ix22302 : mux21_ni port map ( Y=>nx22301, A0=>
      label_9_input_state_machine_3, A1=>data_in(131), S0=>nx42795);
   ix34681 : xor2 port map ( Y=>nx34680, A0=>nx34354, A1=>label_9_output_4);
   ix34685 : xnor2 port map ( Y=>nx34684, A0=>nx34364, A1=>nx34694);
   ix22352 : mux21_ni port map ( Y=>nx22351, A0=>label_9_output_5, A1=>
      label_9_input_5, S0=>nx43521);
   ix5231 : mux21_ni port map ( Y=>nx5230, A0=>nx5226, A1=>
      label_9_input_state_machine_5, S0=>nx43067);
   ix22342 : mux21_ni port map ( Y=>nx22341, A0=>
      label_9_input_state_machine_5, A1=>data_in(133), S0=>nx43361);
   ix34696 : xor2 port map ( Y=>nx34695, A0=>nx34384, A1=>label_9_output_6);
   ix34700 : xnor2 port map ( Y=>nx34699, A0=>nx34403, A1=>nx34709);
   ix22392 : mux21_ni port map ( Y=>nx22391, A0=>label_9_output_7, A1=>
      label_9_input_7, S0=>nx43521);
   ix5295 : mux21_ni port map ( Y=>nx5294, A0=>nx5290, A1=>
      label_9_input_state_machine_7, S0=>nx43067);
   ix22382 : mux21_ni port map ( Y=>nx22381, A0=>
      label_9_input_state_machine_7, A1=>data_in(135), S0=>nx43361);
   ix34711 : xor2 port map ( Y=>nx34710, A0=>nx34436, A1=>label_9_output_8);
   ix34715 : xnor2 port map ( Y=>nx34714, A0=>nx34441, A1=>nx34724);
   ix22432 : mux21_ni port map ( Y=>nx22431, A0=>label_9_output_9, A1=>
      label_9_input_9, S0=>nx43521);
   ix5359 : mux21_ni port map ( Y=>nx5358, A0=>nx5354, A1=>
      label_9_input_state_machine_9, S0=>nx43067);
   ix22422 : mux21_ni port map ( Y=>nx22421, A0=>
      label_9_input_state_machine_9, A1=>data_in(137), S0=>nx43361);
   ix34726 : xor2 port map ( Y=>nx34725, A0=>nx34472, A1=>label_9_output_10
   );
   ix34730 : xnor2 port map ( Y=>nx34729, A0=>nx34477, A1=>nx34739);
   ix22472 : mux21_ni port map ( Y=>nx22471, A0=>label_9_output_11, A1=>
      label_9_input_11, S0=>nx43521);
   ix5423 : mux21_ni port map ( Y=>nx5422, A0=>nx5418, A1=>
      label_9_input_state_machine_11, S0=>nx43069);
   ix22462 : mux21_ni port map ( Y=>nx22461, A0=>
      label_9_input_state_machine_11, A1=>data_in(139), S0=>nx43361);
   ix34741 : xor2 port map ( Y=>nx34740, A0=>nx34508, A1=>label_9_output_12
   );
   ix34745 : xnor2 port map ( Y=>nx34744, A0=>nx34513, A1=>nx34754);
   ix22512 : mux21_ni port map ( Y=>nx22511, A0=>label_9_output_13, A1=>
      label_9_input_13, S0=>nx43521);
   ix5487 : mux21_ni port map ( Y=>nx5486, A0=>nx5482, A1=>
      label_9_input_state_machine_13, S0=>nx43069);
   ix22502 : mux21_ni port map ( Y=>nx22501, A0=>
      label_9_input_state_machine_13, A1=>data_in(141), S0=>nx43361);
   ix34756 : xor2 port map ( Y=>nx34755, A0=>nx34544, A1=>label_9_output_14
   );
   ix5533 : xnor2 port map ( Y=>nx5532, A0=>nx34760, A1=>nx34125);
   ix34770 : xnor2 port map ( Y=>nx34769, A0=>nx34773, A1=>
      max_calc_comparator_fifth_inp1_13);
   ix34776 : or03 port map ( Y=>nx34775, A0=>nx34089, A1=>nx42975, A2=>
      nx42539);
   ix34781 : or03 port map ( Y=>nx34780, A0=>nx34754, A1=>nx42975, A2=>
      nx42539);
   ix5569 : xnor2 port map ( Y=>nx5568, A0=>nx34784, A1=>nx34791);
   ix34798 : xnor2 port map ( Y=>nx34797, A0=>nx34801, A1=>
      max_calc_comparator_fifth_inp1_11);
   ix34804 : or03 port map ( Y=>nx34803, A0=>nx34074, A1=>nx42975, A2=>
      nx42539);
   ix34809 : or03 port map ( Y=>nx34808, A0=>nx34739, A1=>nx42977, A2=>
      nx42539);
   ix5605 : xnor2 port map ( Y=>nx5604, A0=>nx34812, A1=>nx34819);
   ix34826 : xnor2 port map ( Y=>nx34825, A0=>nx34829, A1=>
      max_calc_comparator_fifth_inp1_9);
   ix34832 : or03 port map ( Y=>nx34831, A0=>nx34059, A1=>nx42977, A2=>
      nx43207);
   ix34837 : or03 port map ( Y=>nx34836, A0=>nx34724, A1=>nx42977, A2=>
      nx43207);
   ix5641 : xnor2 port map ( Y=>nx5640, A0=>nx34840, A1=>nx34847);
   ix34854 : xnor2 port map ( Y=>nx34853, A0=>nx34857, A1=>
      max_calc_comparator_fifth_inp1_7);
   ix34860 : or03 port map ( Y=>nx34859, A0=>nx34044, A1=>nx42977, A2=>
      nx43207);
   ix34865 : or03 port map ( Y=>nx34864, A0=>nx34709, A1=>nx42977, A2=>
      nx43207);
   ix5677 : xnor2 port map ( Y=>nx5676, A0=>nx34868, A1=>nx34875);
   ix34882 : xnor2 port map ( Y=>nx34881, A0=>nx34885, A1=>
      max_calc_comparator_fifth_inp1_5);
   ix34888 : or03 port map ( Y=>nx34887, A0=>nx34029, A1=>nx42977, A2=>
      nx43207);
   ix34893 : or03 port map ( Y=>nx34892, A0=>nx34694, A1=>nx42977, A2=>
      nx43207);
   ix5713 : xnor2 port map ( Y=>nx5712, A0=>nx34896, A1=>nx34903);
   ix34910 : xnor2 port map ( Y=>nx34909, A0=>nx34913, A1=>
      max_calc_comparator_fifth_inp1_3);
   ix34916 : or03 port map ( Y=>nx34915, A0=>nx34014, A1=>nx42979, A2=>
      nx43207);
   ix34921 : or03 port map ( Y=>nx34920, A0=>nx34679, A1=>nx42979, A2=>
      nx42541);
   ix5749 : xnor2 port map ( Y=>nx5748, A0=>nx34924, A1=>nx34931);
   ix34942 : or03 port map ( Y=>nx34941, A0=>nx33999, A1=>nx42979, A2=>
      nx42541);
   ix34947 : or03 port map ( Y=>nx34946, A0=>nx34664, A1=>nx42979, A2=>
      nx42541);
   ix5767 : xnor2 port map ( Y=>nx5766, A0=>nx34939, A1=>nx34943);
   ix5977 : xnor2 port map ( Y=>nx5976, A0=>nx34965, A1=>nx34971);
   ix34968 : or03 port map ( Y=>nx34967, A0=>nx34095, A1=>nx42979, A2=>
      nx42541);
   ix34974 : or03 port map ( Y=>nx34973, A0=>nx34987, A1=>nx42979, A2=>
      nx42541);
   ix22852 : mux21_ni port map ( Y=>nx22851, A0=>label_9_output_15, A1=>
      label_9_input_15, S0=>nx43521);
   ix5957 : mux21_ni port map ( Y=>nx5956, A0=>nx5952, A1=>
      label_9_input_state_machine_15, S0=>nx43069);
   ix22842 : mux21_ni port map ( Y=>nx22841, A0=>
      label_9_input_state_machine_15, A1=>data_in(143), S0=>nx43361);
   ix5951 : xnor2 port map ( Y=>nx5950, A0=>nx34549, A1=>label_9_output_15);
   ix34990 : nor04 port map ( Y=>nx2862, A0=>rst, A1=>nx31896, A2=>
      max_calc_state_0, A3=>nx42845);
   ix2857 : oai21 port map ( Y=>nx42845, A0=>nx43453, A1=>max_calc_state_2, 
      B0=>nx42927);
   ix30452 : mux21_ni port map ( Y=>nx30451, A0=>
      max_calc_comparator_first_inp2_14, A1=>nx18156, S0=>nx43391);
   ix18157 : mux21_ni port map ( Y=>nx18156, A0=>nx18152, A1=>nx17622, S0=>
      nx43031);
   ix17623 : mux21_ni port map ( Y=>nx17622, A0=>max_calc_ans2_14, A1=>
      label_2_output_14, S0=>nx43143);
   ix23712 : mux21_ni port map ( Y=>nx23711, A0=>label_2_output_14, A1=>
      label_2_input_14, S0=>nx43413);
   ix7303 : mux21_ni port map ( Y=>nx7302, A0=>nx7298, A1=>
      label_2_input_state_machine_14, S0=>nx43069);
   ix22892 : mux21_ni port map ( Y=>nx22891, A0=>
      label_2_input_state_machine_14, A1=>data_in(30), S0=>nx43361);
   ix23682 : mux21_ni port map ( Y=>nx23681, A0=>label_2_output_12, A1=>
      label_2_input_12, S0=>nx43413);
   ix7245 : mux21_ni port map ( Y=>nx7244, A0=>nx7240, A1=>
      label_2_input_state_machine_12, S0=>nx43069);
   ix23672 : mux21_ni port map ( Y=>nx23671, A0=>
      label_2_input_state_machine_12, A1=>data_in(28), S0=>nx43363);
   ix23642 : mux21_ni port map ( Y=>nx23641, A0=>label_2_output_10, A1=>
      label_2_input_10, S0=>nx43413);
   ix7181 : mux21_ni port map ( Y=>nx7180, A0=>nx7176, A1=>
      label_2_input_state_machine_10, S0=>nx43069);
   ix23632 : mux21_ni port map ( Y=>nx23631, A0=>
      label_2_input_state_machine_10, A1=>data_in(26), S0=>nx43363);
   ix23602 : mux21_ni port map ( Y=>nx23601, A0=>label_2_output_8, A1=>
      label_2_input_8, S0=>nx43413);
   ix7117 : mux21_ni port map ( Y=>nx7116, A0=>nx7112, A1=>
      label_2_input_state_machine_8, S0=>nx43069);
   ix23592 : mux21_ni port map ( Y=>nx23591, A0=>
      label_2_input_state_machine_8, A1=>data_in(24), S0=>nx43363);
   ix23562 : mux21_ni port map ( Y=>nx23561, A0=>label_2_output_6, A1=>
      label_2_input_6, S0=>nx43413);
   ix7053 : mux21_ni port map ( Y=>nx7052, A0=>nx7048, A1=>
      label_2_input_state_machine_6, S0=>nx43071);
   ix23552 : mux21_ni port map ( Y=>nx23551, A0=>
      label_2_input_state_machine_6, A1=>data_in(22), S0=>nx43363);
   ix23522 : mux21_ni port map ( Y=>nx23521, A0=>label_2_output_4, A1=>
      label_2_input_4, S0=>nx43413);
   ix6989 : mux21_ni port map ( Y=>nx6988, A0=>nx6984, A1=>
      label_2_input_state_machine_4, S0=>nx43071);
   ix23512 : mux21_ni port map ( Y=>nx23511, A0=>
      label_2_input_state_machine_4, A1=>data_in(20), S0=>nx43363);
   ix23482 : mux21_ni port map ( Y=>nx23481, A0=>label_2_output_2, A1=>
      label_2_input_2, S0=>nx43413);
   ix6925 : mux21_ni port map ( Y=>nx6924, A0=>nx6920, A1=>
      label_2_input_state_machine_2, S0=>nx43071);
   ix23472 : mux21_ni port map ( Y=>nx23471, A0=>
      label_2_input_state_machine_2, A1=>data_in(18), S0=>nx43363);
   ix23442 : mux21_ni port map ( Y=>nx23441, A0=>label_2_output_0, A1=>
      label_2_input_0, S0=>nx43521);
   ix23432 : mux21_ni port map ( Y=>nx23431, A0=>
      label_2_input_state_machine_0, A1=>data_in(16), S0=>nx43363);
   ix23422 : mux21_ni port map ( Y=>nx23421, A0=>
      booth_booth_integration_output_1_12, A1=>nx6844, S0=>nx43221);
   ix6845 : mux21_ni port map ( Y=>nx6844, A0=>nx41807, A1=>
      booth_booth_integration_output_1_13, S0=>nx43229);
   ix23412 : mux21_ni port map ( Y=>nx23411, A0=>
      booth_booth_integration_output_1_13, A1=>nx6832, S0=>nx43221);
   ix6833 : mux21_ni port map ( Y=>nx6832, A0=>nx41803, A1=>
      booth_booth_integration_output_1_14, S0=>nx43229);
   ix23402 : mux21_ni port map ( Y=>nx23401, A0=>
      booth_booth_integration_output_1_14, A1=>nx6820, S0=>nx43221);
   ix6821 : mux21_ni port map ( Y=>nx6820, A0=>nx41799, A1=>
      booth_booth_integration_output_1_15, S0=>nx43229);
   ix23392 : mux21 port map ( Y=>nx23391, A0=>nx35517, A1=>nx35098, S0=>
      nx43221);
   ix22922 : mux21_ni port map ( Y=>nx22921, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_0, A1=>nx41919, S0=>nx42937
   );
   ix22908 : and02 port map ( Y=>nx22907, A0=>nx43475, A1=>
      booth_booth_integrtaion_1_shift_Reg_count_0);
   ix23102 : mux21_ni port map ( Y=>nx23101, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_9, A1=>nx41905, S0=>nx42937
   );
   ix23092 : mux21_ni port map ( Y=>nx23091, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_9, A1=>output_8_dup_12716, 
      S0=>nx43221);
   ix23082 : mux21_ni port map ( Y=>nx23081, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_8, A1=>output_8_dup_12716, 
      S0=>nx42937);
   ix23072 : mux21_ni port map ( Y=>nx23071, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_8, A1=>output_7_dup_12717, 
      S0=>nx43221);
   ix23062 : mux21_ni port map ( Y=>nx23061, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_7, A1=>output_7_dup_12717, 
      S0=>nx42937);
   ix23052 : mux21_ni port map ( Y=>nx23051, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_7, A1=>output_6_dup_12718, 
      S0=>nx43223);
   ix23042 : mux21_ni port map ( Y=>nx23041, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_6, A1=>output_6_dup_12718, 
      S0=>nx42937);
   ix23032 : mux21_ni port map ( Y=>nx23031, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_6, A1=>output_5_dup_12719, 
      S0=>nx43223);
   ix23022 : mux21_ni port map ( Y=>nx23021, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_5, A1=>output_5_dup_12719, 
      S0=>nx42937);
   ix23012 : mux21_ni port map ( Y=>nx23011, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_5, A1=>output_4_dup_12720, 
      S0=>nx43223);
   ix23002 : mux21_ni port map ( Y=>nx23001, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_4, A1=>output_4_dup_12720, 
      S0=>nx42939);
   ix22992 : mux21_ni port map ( Y=>nx22991, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_4, A1=>output_3_dup_12721, 
      S0=>nx43223);
   ix22982 : mux21_ni port map ( Y=>nx22981, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_3, A1=>output_3_dup_12721, 
      S0=>nx42939);
   ix22972 : mux21_ni port map ( Y=>nx22971, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_3, A1=>output_2_dup_12722, 
      S0=>nx43223);
   ix22962 : mux21_ni port map ( Y=>nx22961, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_2, A1=>output_2_dup_12722, 
      S0=>nx42939);
   ix22952 : mux21_ni port map ( Y=>nx22951, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_2, A1=>output_1_dup_12723, 
      S0=>nx43223);
   ix22942 : mux21_ni port map ( Y=>nx22941, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_1, A1=>output_1_dup_12723, 
      S0=>nx42939);
   ix22932 : mux21_ni port map ( Y=>nx22931, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_1, A1=>nx41919, S0=>nx43223
   );
   ix6261 : nand02 port map ( Y=>nx35244, A0=>nx35171, A1=>
      booth_output_0_dup_12130);
   ix35174 : or03 port map ( Y=>nx35173, A0=>nx35222, A1=>
      booth_booth_integrtaion_1_shift_reg_output_0, A2=>nx43475);
   ix23222 : mux21_ni port map ( Y=>nx23221, A0=>booth_output_0_dup_12130, 
      A1=>nx6240, S0=>nx43225);
   ix6241 : mux21_ni port map ( Y=>nx6240, A0=>nx41781, A1=>
      booth_output_1_dup_12129, S0=>nx43231);
   ix23212 : mux21_ni port map ( Y=>nx23211, A0=>booth_output_1_dup_12129, 
      A1=>nx6228, S0=>nx43225);
   ix6229 : mux21_ni port map ( Y=>nx6228, A0=>nx41777, A1=>
      booth_output_2_dup_12128, S0=>nx43231);
   ix23202 : mux21_ni port map ( Y=>nx23201, A0=>booth_output_2_dup_12128, 
      A1=>nx6216, S0=>nx43225);
   ix6217 : mux21_ni port map ( Y=>nx6216, A0=>nx41773, A1=>
      booth_output_3_dup_12127, S0=>nx43231);
   ix23192 : mux21_ni port map ( Y=>nx23191, A0=>booth_output_3_dup_12127, 
      A1=>nx6204, S0=>nx43225);
   ix6205 : mux21_ni port map ( Y=>nx6204, A0=>nx41769, A1=>
      booth_output_4_dup_12126, S0=>nx43231);
   ix23182 : mux21_ni port map ( Y=>nx23181, A0=>booth_output_4_dup_12126, 
      A1=>nx6192, S0=>nx43225);
   ix6193 : mux21_ni port map ( Y=>nx6192, A0=>nx41765, A1=>
      booth_output_5_dup_12125, S0=>nx43231);
   ix23172 : mux21_ni port map ( Y=>nx23171, A0=>booth_output_5_dup_12125, 
      A1=>nx6180, S0=>nx43225);
   ix6181 : mux21_ni port map ( Y=>nx6180, A0=>nx41761, A1=>
      booth_output_6_dup_12124, S0=>nx43231);
   ix23162 : mux21_ni port map ( Y=>nx23161, A0=>booth_output_6_dup_12124, 
      A1=>nx6168, S0=>nx43225);
   ix6169 : mux21_ni port map ( Y=>nx6168, A0=>nx41757, A1=>
      booth_output_7_dup_12123, S0=>nx43231);
   ix23152 : mux21_ni port map ( Y=>nx23151, A0=>booth_output_7_dup_12123, 
      A1=>nx6156, S0=>nx43227);
   ix6157 : mux21_ni port map ( Y=>nx6156, A0=>nx41753, A1=>
      booth_output_8_dup_12122, S0=>nx43233);
   ix23142 : mux21_ni port map ( Y=>nx23141, A0=>booth_output_8_dup_12122, 
      A1=>nx6144, S0=>nx43227);
   ix6145 : mux21_ni port map ( Y=>nx6144, A0=>nx41749, A1=>
      booth_output_9_dup_12121, S0=>nx43233);
   ix23132 : mux21_ni port map ( Y=>nx23131, A0=>booth_output_9_dup_12121, 
      A1=>nx6132, S0=>nx43227);
   ix6133 : mux21_ni port map ( Y=>nx6132, A0=>nx41745, A1=>
      booth_output_10_dup_12120, S0=>nx43233);
   ix23122 : mux21_ni port map ( Y=>nx23121, A0=>booth_output_10_dup_12120, 
      A1=>nx6120, S0=>nx43227);
   ix6121 : mux21_ni port map ( Y=>nx6120, A0=>nx41741, A1=>
      booth_output_11_dup_12119, S0=>nx43233);
   ix23112 : mux21_ni port map ( Y=>nx23111, A0=>booth_output_11_dup_12119, 
      A1=>nx6108, S0=>nx43227);
   ix6109 : mux21_ni port map ( Y=>nx6108, A0=>nx41729, A1=>
      booth_booth_integration_output_1_12, S0=>nx43233);
   ix23382 : mux21_ni port map ( Y=>nx23381, A0=>
      booth_booth_integration_output_1_16, A1=>nx6790, S0=>nx43227);
   ix6791 : nor02ii port map ( Y=>nx6790, A0=>nx35228, A1=>nx43233);
   ix6267 : nor02ii port map ( Y=>nx6266, A0=>nx35166, A1=>
      booth_booth_integration_output_1_16);
   ix6785 : xor2 port map ( Y=>nx18297, A0=>nx35234, A1=>nx35510);
   ix35250 : or02 port map ( Y=>nx35249, A0=>nx35171, A1=>
      booth_output_0_dup_12130);
   ix6773 : xor2 port map ( Y=>nx18299, A0=>nx35254, A1=>nx42563);
   ix35270 : xor2 port map ( Y=>nx35269, A0=>nx35273, A1=>nx6338);
   ix35282 : nor02ii port map ( Y=>nx35281, A0=>nx6304, A1=>data_in(19));
   ix6749 : xor2 port map ( Y=>nx18301, A0=>nx35306, A1=>nx42565);
   ix23342 : mux21_ni port map ( Y=>nx23341, A0=>
      booth_booth_integration_output_1_20, A1=>nx6742, S0=>nx43227);
   ix6743 : nor02ii port map ( Y=>nx6742, A0=>nx35292, A1=>nx43233);
   ix6737 : xor2 port map ( Y=>nx18302, A0=>nx35311, A1=>nx35507);
   ix6725 : xor2 port map ( Y=>nx18303, A0=>nx35342, A1=>nx42567);
   ix23322 : mux21_ni port map ( Y=>nx23321, A0=>
      booth_booth_integration_output_1_22, A1=>nx6718, S0=>nx42557);
   ix6719 : nor02ii port map ( Y=>nx6718, A0=>nx35328, A1=>nx42561);
   ix6713 : xor2 port map ( Y=>nx18304, A0=>nx35347, A1=>nx35504);
   ix6701 : xor2 port map ( Y=>nx18305, A0=>nx35378, A1=>nx42569);
   ix23302 : mux21_ni port map ( Y=>nx23301, A0=>
      booth_booth_integration_output_1_24, A1=>nx6694, S0=>nx42557);
   ix6695 : nor02ii port map ( Y=>nx6694, A0=>nx35364, A1=>nx42561);
   ix6689 : xor2 port map ( Y=>nx18307, A0=>nx35383, A1=>nx35501);
   ix6677 : xor2 port map ( Y=>nx18309, A0=>nx35414, A1=>nx42571);
   ix23282 : mux21_ni port map ( Y=>nx23281, A0=>
      booth_booth_integration_output_1_26, A1=>nx6670, S0=>nx42557);
   ix6671 : nor02ii port map ( Y=>nx6670, A0=>nx35400, A1=>nx42561);
   ix6665 : xor2 port map ( Y=>nx18311, A0=>nx35419, A1=>nx35498);
   ix6653 : xor2 port map ( Y=>nx18313, A0=>nx35450, A1=>nx42573);
   ix23262 : mux21_ni port map ( Y=>nx23261, A0=>booth_output_28_dup_12118, 
      A1=>nx6646, S0=>nx42557);
   ix6647 : nor02ii port map ( Y=>nx6646, A0=>nx35436, A1=>nx42561);
   ix6641 : xor2 port map ( Y=>nx18315, A0=>nx35455, A1=>nx35495);
   ix6629 : xor2 port map ( Y=>nx18317, A0=>nx35471, A1=>nx42575);
   ix35489 : xor2 port map ( Y=>nx35488, A0=>nx35471, A1=>nx6614);
   ix6803 : nor02ii port map ( Y=>nx6802, A0=>nx6266, A1=>nx42561);
   ix35525 : xnor2 port map ( Y=>nx35524, A0=>nx35520, A1=>nx35534);
   ix23462 : mux21_ni port map ( Y=>nx23461, A0=>label_2_output_1, A1=>
      label_2_input_1, S0=>nx43415);
   ix6893 : mux21_ni port map ( Y=>nx6892, A0=>nx6888, A1=>
      label_2_input_state_machine_1, S0=>nx43071);
   ix23452 : mux21_ni port map ( Y=>nx23451, A0=>
      label_2_input_state_machine_1, A1=>data_in(17), S0=>nx43365);
   ix35540 : xnor2 port map ( Y=>nx35539, A0=>nx35517, A1=>nx35549);
   ix23502 : mux21_ni port map ( Y=>nx23501, A0=>label_2_output_3, A1=>
      label_2_input_3, S0=>nx43415);
   ix6957 : mux21_ni port map ( Y=>nx6956, A0=>nx6952, A1=>
      label_2_input_state_machine_3, S0=>nx43071);
   ix23492 : mux21_ni port map ( Y=>nx23491, A0=>
      label_2_input_state_machine_3, A1=>data_in(19), S0=>nx43365);
   ix35551 : xor2 port map ( Y=>nx35550, A0=>nx35224, A1=>label_2_output_4);
   ix35555 : xnor2 port map ( Y=>nx35554, A0=>nx35234, A1=>nx35564);
   ix23542 : mux21_ni port map ( Y=>nx23541, A0=>label_2_output_5, A1=>
      label_2_input_5, S0=>nx43415);
   ix7021 : mux21_ni port map ( Y=>nx7020, A0=>nx7016, A1=>
      label_2_input_state_machine_5, S0=>nx43071);
   ix23532 : mux21_ni port map ( Y=>nx23531, A0=>
      label_2_input_state_machine_5, A1=>data_in(21), S0=>nx43365);
   ix35566 : xor2 port map ( Y=>nx35565, A0=>nx35254, A1=>label_2_output_6);
   ix35570 : xnor2 port map ( Y=>nx35569, A0=>nx35273, A1=>nx35579);
   ix23582 : mux21_ni port map ( Y=>nx23581, A0=>label_2_output_7, A1=>
      label_2_input_7, S0=>nx43415);
   ix7085 : mux21_ni port map ( Y=>nx7084, A0=>nx7080, A1=>
      label_2_input_state_machine_7, S0=>nx43071);
   ix23572 : mux21_ni port map ( Y=>nx23571, A0=>
      label_2_input_state_machine_7, A1=>data_in(23), S0=>nx43365);
   ix35581 : xor2 port map ( Y=>nx35580, A0=>nx35306, A1=>label_2_output_8);
   ix35585 : xnor2 port map ( Y=>nx35584, A0=>nx35311, A1=>nx35594);
   ix23622 : mux21_ni port map ( Y=>nx23621, A0=>label_2_output_9, A1=>
      label_2_input_9, S0=>nx43415);
   ix7149 : mux21_ni port map ( Y=>nx7148, A0=>nx7144, A1=>
      label_2_input_state_machine_9, S0=>nx42289);
   ix23612 : mux21_ni port map ( Y=>nx23611, A0=>
      label_2_input_state_machine_9, A1=>data_in(25), S0=>nx43365);
   ix35596 : xor2 port map ( Y=>nx35595, A0=>nx35342, A1=>label_2_output_10
   );
   ix35600 : xnor2 port map ( Y=>nx35599, A0=>nx35347, A1=>nx35609);
   ix23662 : mux21_ni port map ( Y=>nx23661, A0=>label_2_output_11, A1=>
      label_2_input_11, S0=>nx43415);
   ix7213 : mux21_ni port map ( Y=>nx7212, A0=>nx7208, A1=>
      label_2_input_state_machine_11, S0=>nx42289);
   ix23652 : mux21_ni port map ( Y=>nx23651, A0=>
      label_2_input_state_machine_11, A1=>data_in(27), S0=>nx43365);
   ix35611 : xor2 port map ( Y=>nx35610, A0=>nx35378, A1=>label_2_output_12
   );
   ix35615 : xnor2 port map ( Y=>nx35614, A0=>nx35383, A1=>nx35624);
   ix23702 : mux21_ni port map ( Y=>nx23701, A0=>label_2_output_13, A1=>
      label_2_input_13, S0=>nx43415);
   ix7277 : mux21_ni port map ( Y=>nx7276, A0=>nx7272, A1=>
      label_2_input_state_machine_13, S0=>nx42289);
   ix23692 : mux21_ni port map ( Y=>nx23691, A0=>
      label_2_input_state_machine_13, A1=>data_in(29), S0=>nx43365);
   ix35626 : xor2 port map ( Y=>nx35625, A0=>nx35414, A1=>label_2_output_14
   );
   ix30102 : mux21_ni port map ( Y=>nx30101, A0=>nx17612, A1=>
      max_calc_ans2_14, S0=>nx42991);
   ix17613 : mux21 port map ( Y=>nx17612, A0=>nx37785, A1=>nx35633, S0=>
      nx43019);
   ix11809 : mux21_ni port map ( Y=>nx11808, A0=>max_calc_ans3_14, A1=>
      label_3_output_14, S0=>nx43137);
   ix24542 : mux21_ni port map ( Y=>nx24541, A0=>label_3_output_14, A1=>
      label_3_input_14, S0=>nx43417);
   ix8613 : mux21_ni port map ( Y=>nx8612, A0=>nx8608, A1=>
      label_3_input_state_machine_14, S0=>nx43073);
   ix23722 : mux21_ni port map ( Y=>nx23721, A0=>
      label_3_input_state_machine_14, A1=>data_in(46), S0=>nx43367);
   ix24512 : mux21_ni port map ( Y=>nx24511, A0=>label_3_output_12, A1=>
      label_3_input_12, S0=>nx43417);
   ix8555 : mux21_ni port map ( Y=>nx8554, A0=>nx8550, A1=>
      label_3_input_state_machine_12, S0=>nx43073);
   ix24502 : mux21_ni port map ( Y=>nx24501, A0=>
      label_3_input_state_machine_12, A1=>data_in(44), S0=>nx43367);
   ix24472 : mux21_ni port map ( Y=>nx24471, A0=>label_3_output_10, A1=>
      label_3_input_10, S0=>nx43417);
   ix8491 : mux21_ni port map ( Y=>nx8490, A0=>nx8486, A1=>
      label_3_input_state_machine_10, S0=>nx43073);
   ix24462 : mux21_ni port map ( Y=>nx24461, A0=>
      label_3_input_state_machine_10, A1=>data_in(42), S0=>nx43367);
   ix24432 : mux21_ni port map ( Y=>nx24431, A0=>label_3_output_8, A1=>
      label_3_input_8, S0=>nx43417);
   ix8427 : mux21_ni port map ( Y=>nx8426, A0=>nx8422, A1=>
      label_3_input_state_machine_8, S0=>nx43073);
   ix24422 : mux21_ni port map ( Y=>nx24421, A0=>
      label_3_input_state_machine_8, A1=>data_in(40), S0=>nx43367);
   ix24392 : mux21_ni port map ( Y=>nx24391, A0=>label_3_output_6, A1=>
      label_3_input_6, S0=>nx43417);
   ix8363 : mux21_ni port map ( Y=>nx8362, A0=>nx8358, A1=>
      label_3_input_state_machine_6, S0=>nx43075);
   ix24382 : mux21_ni port map ( Y=>nx24381, A0=>
      label_3_input_state_machine_6, A1=>data_in(38), S0=>nx43367);
   ix24352 : mux21_ni port map ( Y=>nx24351, A0=>label_3_output_4, A1=>
      label_3_input_4, S0=>nx43417);
   ix8299 : mux21_ni port map ( Y=>nx8298, A0=>nx8294, A1=>
      label_3_input_state_machine_4, S0=>nx42289);
   ix24342 : mux21_ni port map ( Y=>nx24341, A0=>
      label_3_input_state_machine_4, A1=>data_in(36), S0=>nx43367);
   ix24312 : mux21_ni port map ( Y=>nx24311, A0=>label_3_output_2, A1=>
      label_3_input_2, S0=>nx43417);
   ix8235 : mux21_ni port map ( Y=>nx8234, A0=>nx8230, A1=>
      label_3_input_state_machine_2, S0=>nx42289);
   ix24302 : mux21_ni port map ( Y=>nx24301, A0=>
      label_3_input_state_machine_2, A1=>data_in(34), S0=>nx43367);
   ix24272 : mux21_ni port map ( Y=>nx24271, A0=>label_3_output_0, A1=>
      label_3_input_0, S0=>nx43419);
   ix24262 : mux21_ni port map ( Y=>nx24261, A0=>
      label_3_input_state_machine_0, A1=>data_in(32), S0=>nx43369);
   ix24252 : mux21_ni port map ( Y=>nx24251, A0=>
      booth_booth_integration_output_2_12, A1=>nx8154, S0=>nx43235);
   ix8155 : mux21_ni port map ( Y=>nx8154, A0=>nx41807, A1=>
      booth_booth_integration_output_2_13, S0=>nx43243);
   ix24242 : mux21_ni port map ( Y=>nx24241, A0=>
      booth_booth_integration_output_2_13, A1=>nx8142, S0=>nx43235);
   ix8143 : mux21_ni port map ( Y=>nx8142, A0=>nx41803, A1=>
      booth_booth_integration_output_2_14, S0=>nx43243);
   ix24232 : mux21_ni port map ( Y=>nx24231, A0=>
      booth_booth_integration_output_2_14, A1=>nx8130, S0=>nx43235);
   ix8131 : mux21_ni port map ( Y=>nx8130, A0=>nx41799, A1=>
      booth_booth_integration_output_2_15, S0=>nx43243);
   ix24222 : mux21 port map ( Y=>nx24221, A0=>nx36155, A1=>nx35736, S0=>
      nx43235);
   ix23752 : mux21_ni port map ( Y=>nx23751, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_0, A1=>nx41951, S0=>nx42941
   );
   ix23738 : and02 port map ( Y=>nx23737, A0=>nx43479, A1=>
      booth_booth_integrtaion_2_shift_Reg_count_0);
   ix23932 : mux21_ni port map ( Y=>nx23931, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_9, A1=>nx41937, S0=>nx42941
   );
   ix23922 : mux21_ni port map ( Y=>nx23921, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_9, A1=>output_8_dup_12744, 
      S0=>nx43235);
   ix23912 : mux21_ni port map ( Y=>nx23911, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_8, A1=>output_8_dup_12744, 
      S0=>nx42941);
   ix23902 : mux21_ni port map ( Y=>nx23901, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_8, A1=>output_7_dup_12745, 
      S0=>nx43235);
   ix23892 : mux21_ni port map ( Y=>nx23891, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_7, A1=>output_7_dup_12745, 
      S0=>nx42941);
   ix23882 : mux21_ni port map ( Y=>nx23881, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_7, A1=>output_6_dup_12746, 
      S0=>nx43237);
   ix23872 : mux21_ni port map ( Y=>nx23871, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_6, A1=>output_6_dup_12746, 
      S0=>nx42941);
   ix23862 : mux21_ni port map ( Y=>nx23861, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_6, A1=>output_5_dup_12747, 
      S0=>nx43237);
   ix23852 : mux21_ni port map ( Y=>nx23851, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_5, A1=>output_5_dup_12747, 
      S0=>nx42941);
   ix23842 : mux21_ni port map ( Y=>nx23841, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_5, A1=>output_4_dup_12748, 
      S0=>nx43237);
   ix23832 : mux21_ni port map ( Y=>nx23831, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_4, A1=>output_4_dup_12748, 
      S0=>nx42943);
   ix23822 : mux21_ni port map ( Y=>nx23821, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_4, A1=>output_3_dup_12749, 
      S0=>nx43237);
   ix23812 : mux21_ni port map ( Y=>nx23811, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_3, A1=>output_3_dup_12749, 
      S0=>nx42943);
   ix23802 : mux21_ni port map ( Y=>nx23801, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_3, A1=>output_2_dup_12750, 
      S0=>nx43237);
   ix23792 : mux21_ni port map ( Y=>nx23791, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_2, A1=>output_2_dup_12750, 
      S0=>nx42943);
   ix23782 : mux21_ni port map ( Y=>nx23781, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_2, A1=>output_1_dup_12751, 
      S0=>nx43237);
   ix23772 : mux21_ni port map ( Y=>nx23771, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_1, A1=>output_1_dup_12751, 
      S0=>nx42943);
   ix23762 : mux21_ni port map ( Y=>nx23761, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_1, A1=>nx41951, S0=>nx43237
   );
   ix7571 : nand02 port map ( Y=>nx35882, A0=>nx35809, A1=>
      booth_output_0_dup_12149);
   ix35812 : or03 port map ( Y=>nx35811, A0=>nx35860, A1=>
      booth_booth_integrtaion_2_shift_reg_output_0, A2=>nx43479);
   ix24052 : mux21_ni port map ( Y=>nx24051, A0=>booth_output_0_dup_12149, 
      A1=>nx7550, S0=>nx43239);
   ix7551 : mux21_ni port map ( Y=>nx7550, A0=>nx41781, A1=>
      booth_output_1_dup_12148, S0=>nx43245);
   ix24042 : mux21_ni port map ( Y=>nx24041, A0=>booth_output_1_dup_12148, 
      A1=>nx7538, S0=>nx43239);
   ix7539 : mux21_ni port map ( Y=>nx7538, A0=>nx41777, A1=>
      booth_output_2_dup_12147, S0=>nx43245);
   ix24032 : mux21_ni port map ( Y=>nx24031, A0=>booth_output_2_dup_12147, 
      A1=>nx7526, S0=>nx43239);
   ix7527 : mux21_ni port map ( Y=>nx7526, A0=>nx41773, A1=>
      booth_output_3_dup_12146, S0=>nx43245);
   ix24022 : mux21_ni port map ( Y=>nx24021, A0=>booth_output_3_dup_12146, 
      A1=>nx7514, S0=>nx43239);
   ix7515 : mux21_ni port map ( Y=>nx7514, A0=>nx41769, A1=>
      booth_output_4_dup_12145, S0=>nx43245);
   ix24012 : mux21_ni port map ( Y=>nx24011, A0=>booth_output_4_dup_12145, 
      A1=>nx7502, S0=>nx43239);
   ix7503 : mux21_ni port map ( Y=>nx7502, A0=>nx41765, A1=>
      booth_output_5_dup_12144, S0=>nx43245);
   ix24002 : mux21_ni port map ( Y=>nx24001, A0=>booth_output_5_dup_12144, 
      A1=>nx7490, S0=>nx43239);
   ix7491 : mux21_ni port map ( Y=>nx7490, A0=>nx41761, A1=>
      booth_output_6_dup_12143, S0=>nx43245);
   ix23992 : mux21_ni port map ( Y=>nx23991, A0=>booth_output_6_dup_12143, 
      A1=>nx7478, S0=>nx43239);
   ix7479 : mux21_ni port map ( Y=>nx7478, A0=>nx41757, A1=>
      booth_output_7_dup_12142, S0=>nx43245);
   ix23982 : mux21_ni port map ( Y=>nx23981, A0=>booth_output_7_dup_12142, 
      A1=>nx7466, S0=>nx43241);
   ix7467 : mux21_ni port map ( Y=>nx7466, A0=>nx41753, A1=>
      booth_output_8_dup_12141, S0=>nx43247);
   ix23972 : mux21_ni port map ( Y=>nx23971, A0=>booth_output_8_dup_12141, 
      A1=>nx7454, S0=>nx43241);
   ix7455 : mux21_ni port map ( Y=>nx7454, A0=>nx41749, A1=>
      booth_output_9_dup_12140, S0=>nx43247);
   ix23962 : mux21_ni port map ( Y=>nx23961, A0=>booth_output_9_dup_12140, 
      A1=>nx7442, S0=>nx43241);
   ix7443 : mux21_ni port map ( Y=>nx7442, A0=>nx41745, A1=>
      booth_output_10_dup_12139, S0=>nx43247);
   ix23952 : mux21_ni port map ( Y=>nx23951, A0=>booth_output_10_dup_12139, 
      A1=>nx7430, S0=>nx43241);
   ix7431 : mux21_ni port map ( Y=>nx7430, A0=>nx41741, A1=>
      booth_output_11_dup_12138, S0=>nx43247);
   ix23942 : mux21_ni port map ( Y=>nx23941, A0=>booth_output_11_dup_12138, 
      A1=>nx7418, S0=>nx43241);
   ix7419 : mux21_ni port map ( Y=>nx7418, A0=>nx41729, A1=>
      booth_booth_integration_output_2_12, S0=>nx43247);
   ix24212 : mux21_ni port map ( Y=>nx24211, A0=>
      booth_booth_integration_output_2_16, A1=>nx8100, S0=>nx43241);
   ix8101 : nor02ii port map ( Y=>nx8100, A0=>nx35866, A1=>nx43247);
   ix7577 : nor02ii port map ( Y=>nx7576, A0=>nx35804, A1=>
      booth_booth_integration_output_2_16);
   ix8095 : xor2 port map ( Y=>nx18337, A0=>nx35872, A1=>nx36148);
   ix35888 : or02 port map ( Y=>nx35887, A0=>nx35809, A1=>
      booth_output_0_dup_12149);
   ix8083 : xor2 port map ( Y=>nx18339, A0=>nx35892, A1=>nx42589);
   ix35908 : xor2 port map ( Y=>nx35907, A0=>nx35911, A1=>nx7648);
   ix35920 : nor02ii port map ( Y=>nx35919, A0=>nx7614, A1=>data_in(35));
   ix8059 : xor2 port map ( Y=>nx18343, A0=>nx35944, A1=>nx42591);
   ix24172 : mux21_ni port map ( Y=>nx24171, A0=>
      booth_booth_integration_output_2_20, A1=>nx8052, S0=>nx43241);
   ix8053 : nor02ii port map ( Y=>nx8052, A0=>nx35930, A1=>nx43247);
   ix8047 : xor2 port map ( Y=>nx18345, A0=>nx35949, A1=>nx36145);
   ix8035 : xor2 port map ( Y=>nx18347, A0=>nx35980, A1=>nx42593);
   ix24152 : mux21_ni port map ( Y=>nx24151, A0=>
      booth_booth_integration_output_2_22, A1=>nx8028, S0=>nx42583);
   ix8029 : nor02ii port map ( Y=>nx8028, A0=>nx35966, A1=>nx42587);
   ix8023 : xor2 port map ( Y=>nx18349, A0=>nx35985, A1=>nx36142);
   ix8011 : xor2 port map ( Y=>nx18350, A0=>nx36016, A1=>nx42595);
   ix24132 : mux21_ni port map ( Y=>nx24131, A0=>
      booth_booth_integration_output_2_24, A1=>nx8004, S0=>nx42583);
   ix8005 : nor02ii port map ( Y=>nx8004, A0=>nx36002, A1=>nx42587);
   ix7999 : xor2 port map ( Y=>nx18351, A0=>nx36021, A1=>nx36139);
   ix7987 : xor2 port map ( Y=>nx18352, A0=>nx36052, A1=>nx42597);
   ix24112 : mux21_ni port map ( Y=>nx24111, A0=>
      booth_booth_integration_output_2_26, A1=>nx7980, S0=>nx42583);
   ix7981 : nor02ii port map ( Y=>nx7980, A0=>nx36038, A1=>nx42587);
   ix7975 : xor2 port map ( Y=>nx18353, A0=>nx36057, A1=>nx36136);
   ix7963 : xor2 port map ( Y=>nx18354, A0=>nx36088, A1=>nx42599);
   ix24092 : mux21_ni port map ( Y=>nx24091, A0=>booth_output_28_dup_12137, 
      A1=>nx7956, S0=>nx42583);
   ix7957 : nor02ii port map ( Y=>nx7956, A0=>nx36074, A1=>nx42587);
   ix7951 : xor2 port map ( Y=>nx18355, A0=>nx36093, A1=>nx36133);
   ix7939 : xor2 port map ( Y=>nx18357, A0=>nx36109, A1=>nx42601);
   ix36127 : xor2 port map ( Y=>nx36126, A0=>nx36109, A1=>nx7924);
   ix8113 : nor02ii port map ( Y=>nx8112, A0=>nx7576, A1=>nx42587);
   ix36163 : xnor2 port map ( Y=>nx36162, A0=>nx36158, A1=>nx36172);
   ix24292 : mux21_ni port map ( Y=>nx24291, A0=>label_3_output_1, A1=>
      label_3_input_1, S0=>nx43419);
   ix8203 : mux21_ni port map ( Y=>nx8202, A0=>nx8198, A1=>
      label_3_input_state_machine_1, S0=>nx42289);
   ix24282 : mux21_ni port map ( Y=>nx24281, A0=>
      label_3_input_state_machine_1, A1=>data_in(33), S0=>nx43369);
   ix36178 : xnor2 port map ( Y=>nx36177, A0=>nx36155, A1=>nx36187);
   ix24332 : mux21_ni port map ( Y=>nx24331, A0=>label_3_output_3, A1=>
      label_3_input_3, S0=>nx43419);
   ix8267 : mux21_ni port map ( Y=>nx8266, A0=>nx8262, A1=>
      label_3_input_state_machine_3, S0=>nx42289);
   ix24322 : mux21_ni port map ( Y=>nx24321, A0=>
      label_3_input_state_machine_3, A1=>data_in(35), S0=>nx43369);
   ix36189 : xor2 port map ( Y=>nx36188, A0=>nx35862, A1=>label_3_output_4);
   ix36193 : xnor2 port map ( Y=>nx36192, A0=>nx35872, A1=>nx36202);
   ix24372 : mux21_ni port map ( Y=>nx24371, A0=>label_3_output_5, A1=>
      label_3_input_5, S0=>nx43419);
   ix8331 : mux21_ni port map ( Y=>nx8330, A0=>nx8326, A1=>
      label_3_input_state_machine_5, S0=>nx43075);
   ix24362 : mux21_ni port map ( Y=>nx24361, A0=>
      label_3_input_state_machine_5, A1=>data_in(37), S0=>nx43369);
   ix36204 : xor2 port map ( Y=>nx36203, A0=>nx35892, A1=>label_3_output_6);
   ix36208 : xnor2 port map ( Y=>nx36207, A0=>nx35911, A1=>nx36217);
   ix24412 : mux21_ni port map ( Y=>nx24411, A0=>label_3_output_7, A1=>
      label_3_input_7, S0=>nx43419);
   ix8395 : mux21_ni port map ( Y=>nx8394, A0=>nx8390, A1=>
      label_3_input_state_machine_7, S0=>nx43075);
   ix24402 : mux21_ni port map ( Y=>nx24401, A0=>
      label_3_input_state_machine_7, A1=>data_in(39), S0=>nx43369);
   ix36219 : xor2 port map ( Y=>nx36218, A0=>nx35944, A1=>label_3_output_8);
   ix36223 : xnor2 port map ( Y=>nx36222, A0=>nx35949, A1=>nx36232);
   ix24452 : mux21_ni port map ( Y=>nx24451, A0=>label_3_output_9, A1=>
      label_3_input_9, S0=>nx43419);
   ix8459 : mux21_ni port map ( Y=>nx8458, A0=>nx8454, A1=>
      label_3_input_state_machine_9, S0=>nx43075);
   ix24442 : mux21_ni port map ( Y=>nx24441, A0=>
      label_3_input_state_machine_9, A1=>data_in(41), S0=>nx43369);
   ix36234 : xor2 port map ( Y=>nx36233, A0=>nx35980, A1=>label_3_output_10
   );
   ix36238 : xnor2 port map ( Y=>nx36237, A0=>nx35985, A1=>nx36247);
   ix24492 : mux21_ni port map ( Y=>nx24491, A0=>label_3_output_11, A1=>
      label_3_input_11, S0=>nx43419);
   ix8523 : mux21_ni port map ( Y=>nx8522, A0=>nx8518, A1=>
      label_3_input_state_machine_11, S0=>nx43075);
   ix24482 : mux21_ni port map ( Y=>nx24481, A0=>
      label_3_input_state_machine_11, A1=>data_in(43), S0=>nx43369);
   ix36249 : xor2 port map ( Y=>nx36248, A0=>nx36016, A1=>label_3_output_12
   );
   ix36253 : xnor2 port map ( Y=>nx36252, A0=>nx36021, A1=>nx36262);
   ix24532 : mux21_ni port map ( Y=>nx24531, A0=>label_3_output_13, A1=>
      label_3_input_13, S0=>nx43421);
   ix8587 : mux21_ni port map ( Y=>nx8586, A0=>nx8582, A1=>
      label_3_input_state_machine_13, S0=>nx43075);
   ix24522 : mux21_ni port map ( Y=>nx24521, A0=>
      label_3_input_state_machine_13, A1=>data_in(45), S0=>nx43371);
   ix36264 : xor2 port map ( Y=>nx36263, A0=>nx36052, A1=>label_3_output_14
   );
   ix11795 : mux21 port map ( Y=>nx11794, A0=>nx36907, A1=>nx36271, S0=>
      nx43007);
   ix25372 : mux21_ni port map ( Y=>nx25371, A0=>label_5_output_14, A1=>
      label_5_input_14, S0=>nx43421);
   ix9933 : mux21_ni port map ( Y=>nx9932, A0=>nx9928, A1=>
      label_5_input_state_machine_14, S0=>nx43075);
   ix24552 : mux21_ni port map ( Y=>nx24551, A0=>
      label_5_input_state_machine_14, A1=>data_in(78), S0=>nx43371);
   ix25342 : mux21_ni port map ( Y=>nx25341, A0=>label_5_output_12, A1=>
      label_5_input_12, S0=>nx43421);
   ix9875 : mux21_ni port map ( Y=>nx9874, A0=>nx9870, A1=>
      label_5_input_state_machine_12, S0=>nx43077);
   ix25332 : mux21_ni port map ( Y=>nx25331, A0=>
      label_5_input_state_machine_12, A1=>data_in(76), S0=>nx43371);
   ix25302 : mux21_ni port map ( Y=>nx25301, A0=>label_5_output_10, A1=>
      label_5_input_10, S0=>nx43421);
   ix9811 : mux21_ni port map ( Y=>nx9810, A0=>nx9806, A1=>
      label_5_input_state_machine_10, S0=>nx43077);
   ix25292 : mux21_ni port map ( Y=>nx25291, A0=>
      label_5_input_state_machine_10, A1=>data_in(74), S0=>nx43371);
   ix25262 : mux21_ni port map ( Y=>nx25261, A0=>label_5_output_8, A1=>
      label_5_input_8, S0=>nx43421);
   ix9747 : mux21_ni port map ( Y=>nx9746, A0=>nx9742, A1=>
      label_5_input_state_machine_8, S0=>nx43077);
   ix25252 : mux21_ni port map ( Y=>nx25251, A0=>
      label_5_input_state_machine_8, A1=>data_in(72), S0=>nx43371);
   ix25222 : mux21_ni port map ( Y=>nx25221, A0=>label_5_output_6, A1=>
      label_5_input_6, S0=>nx43421);
   ix9683 : mux21_ni port map ( Y=>nx9682, A0=>nx9678, A1=>
      label_5_input_state_machine_6, S0=>nx43077);
   ix25212 : mux21_ni port map ( Y=>nx25211, A0=>
      label_5_input_state_machine_6, A1=>data_in(70), S0=>nx43371);
   ix25182 : mux21_ni port map ( Y=>nx25181, A0=>label_5_output_4, A1=>
      label_5_input_4, S0=>nx43421);
   ix9619 : mux21_ni port map ( Y=>nx9618, A0=>nx9614, A1=>
      label_5_input_state_machine_4, S0=>nx43077);
   ix25172 : mux21_ni port map ( Y=>nx25171, A0=>
      label_5_input_state_machine_4, A1=>data_in(68), S0=>nx43371);
   ix25142 : mux21_ni port map ( Y=>nx25141, A0=>label_5_output_2, A1=>
      label_5_input_2, S0=>nx43423);
   ix9555 : mux21_ni port map ( Y=>nx9554, A0=>nx9550, A1=>
      label_5_input_state_machine_2, S0=>nx43077);
   ix25132 : mux21_ni port map ( Y=>nx25131, A0=>
      label_5_input_state_machine_2, A1=>data_in(66), S0=>nx42797);
   ix25102 : mux21_ni port map ( Y=>nx25101, A0=>label_5_output_0, A1=>
      label_5_input_0, S0=>nx43423);
   ix25092 : mux21_ni port map ( Y=>nx25091, A0=>
      label_5_input_state_machine_0, A1=>data_in(64), S0=>nx42797);
   ix25082 : mux21_ni port map ( Y=>nx25081, A0=>
      booth_booth_integration_output_4_12, A1=>nx9474, S0=>nx43249);
   ix9475 : mux21_ni port map ( Y=>nx9474, A0=>nx41807, A1=>
      booth_booth_integration_output_4_13, S0=>nx43257);
   ix25072 : mux21_ni port map ( Y=>nx25071, A0=>
      booth_booth_integration_output_4_13, A1=>nx9462, S0=>nx43249);
   ix9463 : mux21_ni port map ( Y=>nx9462, A0=>nx41803, A1=>
      booth_booth_integration_output_4_14, S0=>nx43257);
   ix25062 : mux21_ni port map ( Y=>nx25061, A0=>
      booth_booth_integration_output_4_14, A1=>nx9450, S0=>nx43249);
   ix9451 : mux21_ni port map ( Y=>nx9450, A0=>nx41799, A1=>
      booth_booth_integration_output_4_15, S0=>nx43257);
   ix25052 : mux21 port map ( Y=>nx25051, A0=>nx36792, A1=>nx36373, S0=>
      nx43249);
   ix24582 : mux21_ni port map ( Y=>nx24581, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_0, A1=>nx41983, S0=>nx42945
   );
   ix24568 : and02 port map ( Y=>nx24567, A0=>nx43483, A1=>
      booth_booth_integrtaion_4_shift_Reg_count_0);
   ix24762 : mux21_ni port map ( Y=>nx24761, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_9, A1=>nx41969, S0=>nx42945
   );
   ix24752 : mux21_ni port map ( Y=>nx24751, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_9, A1=>output_8_dup_12800, 
      S0=>nx43249);
   ix24742 : mux21_ni port map ( Y=>nx24741, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_8, A1=>output_8_dup_12800, 
      S0=>nx42945);
   ix24732 : mux21_ni port map ( Y=>nx24731, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_8, A1=>output_7_dup_12801, 
      S0=>nx43249);
   ix24722 : mux21_ni port map ( Y=>nx24721, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_7, A1=>output_7_dup_12801, 
      S0=>nx42945);
   ix24712 : mux21_ni port map ( Y=>nx24711, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_7, A1=>output_6_dup_12802, 
      S0=>nx43251);
   ix24702 : mux21_ni port map ( Y=>nx24701, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_6, A1=>output_6_dup_12802, 
      S0=>nx42945);
   ix24692 : mux21_ni port map ( Y=>nx24691, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_6, A1=>output_5_dup_12803, 
      S0=>nx43251);
   ix24682 : mux21_ni port map ( Y=>nx24681, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_5, A1=>output_5_dup_12803, 
      S0=>nx42945);
   ix24672 : mux21_ni port map ( Y=>nx24671, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_5, A1=>output_4_dup_12804, 
      S0=>nx43251);
   ix24662 : mux21_ni port map ( Y=>nx24661, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_4, A1=>output_4_dup_12804, 
      S0=>nx42947);
   ix24652 : mux21_ni port map ( Y=>nx24651, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_4, A1=>output_3_dup_12805, 
      S0=>nx43251);
   ix24642 : mux21_ni port map ( Y=>nx24641, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_3, A1=>output_3_dup_12805, 
      S0=>nx42947);
   ix24632 : mux21_ni port map ( Y=>nx24631, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_3, A1=>output_2_dup_12806, 
      S0=>nx43251);
   ix24622 : mux21_ni port map ( Y=>nx24621, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_2, A1=>output_2_dup_12806, 
      S0=>nx42947);
   ix24612 : mux21_ni port map ( Y=>nx24611, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_2, A1=>output_1_dup_12807, 
      S0=>nx43251);
   ix24602 : mux21_ni port map ( Y=>nx24601, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_1, A1=>output_1_dup_12807, 
      S0=>nx42947);
   ix24592 : mux21_ni port map ( Y=>nx24591, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_1, A1=>nx41983, S0=>nx43251
   );
   ix8891 : nand02 port map ( Y=>nx36519, A0=>nx36446, A1=>
      booth_output_0_dup_12187);
   ix36449 : or03 port map ( Y=>nx36448, A0=>nx36497, A1=>
      booth_booth_integrtaion_4_shift_reg_output_0, A2=>nx43483);
   ix24882 : mux21_ni port map ( Y=>nx24881, A0=>booth_output_0_dup_12187, 
      A1=>nx8870, S0=>nx43253);
   ix8871 : mux21_ni port map ( Y=>nx8870, A0=>nx41781, A1=>
      booth_output_1_dup_12186, S0=>nx43259);
   ix24872 : mux21_ni port map ( Y=>nx24871, A0=>booth_output_1_dup_12186, 
      A1=>nx8858, S0=>nx43253);
   ix8859 : mux21_ni port map ( Y=>nx8858, A0=>nx41777, A1=>
      booth_output_2_dup_12185, S0=>nx43259);
   ix24862 : mux21_ni port map ( Y=>nx24861, A0=>booth_output_2_dup_12185, 
      A1=>nx8846, S0=>nx43253);
   ix8847 : mux21_ni port map ( Y=>nx8846, A0=>nx41773, A1=>
      booth_output_3_dup_12184, S0=>nx43259);
   ix24852 : mux21_ni port map ( Y=>nx24851, A0=>booth_output_3_dup_12184, 
      A1=>nx8834, S0=>nx43253);
   ix8835 : mux21_ni port map ( Y=>nx8834, A0=>nx41769, A1=>
      booth_output_4_dup_12183, S0=>nx43259);
   ix24842 : mux21_ni port map ( Y=>nx24841, A0=>booth_output_4_dup_12183, 
      A1=>nx8822, S0=>nx43253);
   ix8823 : mux21_ni port map ( Y=>nx8822, A0=>nx41765, A1=>
      booth_output_5_dup_12182, S0=>nx43259);
   ix24832 : mux21_ni port map ( Y=>nx24831, A0=>booth_output_5_dup_12182, 
      A1=>nx8810, S0=>nx43253);
   ix8811 : mux21_ni port map ( Y=>nx8810, A0=>nx41761, A1=>
      booth_output_6_dup_12181, S0=>nx43259);
   ix24822 : mux21_ni port map ( Y=>nx24821, A0=>booth_output_6_dup_12181, 
      A1=>nx8798, S0=>nx43253);
   ix8799 : mux21_ni port map ( Y=>nx8798, A0=>nx41757, A1=>
      booth_output_7_dup_12180, S0=>nx43259);
   ix24812 : mux21_ni port map ( Y=>nx24811, A0=>booth_output_7_dup_12180, 
      A1=>nx8786, S0=>nx43255);
   ix8787 : mux21_ni port map ( Y=>nx8786, A0=>nx41753, A1=>
      booth_output_8_dup_12179, S0=>nx43261);
   ix24802 : mux21_ni port map ( Y=>nx24801, A0=>booth_output_8_dup_12179, 
      A1=>nx8774, S0=>nx43255);
   ix8775 : mux21_ni port map ( Y=>nx8774, A0=>nx41749, A1=>
      booth_output_9_dup_12178, S0=>nx43261);
   ix24792 : mux21_ni port map ( Y=>nx24791, A0=>booth_output_9_dup_12178, 
      A1=>nx8762, S0=>nx43255);
   ix8763 : mux21_ni port map ( Y=>nx8762, A0=>nx41745, A1=>
      booth_output_10_dup_12177, S0=>nx43261);
   ix24782 : mux21_ni port map ( Y=>nx24781, A0=>booth_output_10_dup_12177, 
      A1=>nx8750, S0=>nx43255);
   ix8751 : mux21_ni port map ( Y=>nx8750, A0=>nx41741, A1=>
      booth_output_11_dup_12176, S0=>nx43261);
   ix24772 : mux21_ni port map ( Y=>nx24771, A0=>booth_output_11_dup_12176, 
      A1=>nx8738, S0=>nx43255);
   ix8739 : mux21_ni port map ( Y=>nx8738, A0=>nx41729, A1=>
      booth_booth_integration_output_4_12, S0=>nx43261);
   ix25042 : mux21_ni port map ( Y=>nx25041, A0=>
      booth_booth_integration_output_4_16, A1=>nx9420, S0=>nx43255);
   ix9421 : nor02ii port map ( Y=>nx9420, A0=>nx36503, A1=>nx43261);
   ix8897 : nor02ii port map ( Y=>nx8896, A0=>nx36441, A1=>
      booth_booth_integration_output_4_16);
   ix9415 : xor2 port map ( Y=>nx18379, A0=>nx36509, A1=>nx36785);
   ix36525 : or02 port map ( Y=>nx36524, A0=>nx36446, A1=>
      booth_output_0_dup_12187);
   ix9403 : xor2 port map ( Y=>nx18380, A0=>nx36529, A1=>nx42615);
   ix36545 : xor2 port map ( Y=>nx36544, A0=>nx36548, A1=>nx8968);
   ix36557 : nor02ii port map ( Y=>nx36556, A0=>nx8934, A1=>data_in(67));
   ix9379 : xor2 port map ( Y=>nx18382, A0=>nx36581, A1=>nx42617);
   ix25002 : mux21_ni port map ( Y=>nx25001, A0=>
      booth_booth_integration_output_4_20, A1=>nx9372, S0=>nx43255);
   ix9373 : nor02ii port map ( Y=>nx9372, A0=>nx36567, A1=>nx43261);
   ix9367 : xor2 port map ( Y=>nx18383, A0=>nx36586, A1=>nx36782);
   ix9355 : xor2 port map ( Y=>nx18385, A0=>nx36617, A1=>nx42619);
   ix24982 : mux21_ni port map ( Y=>nx24981, A0=>
      booth_booth_integration_output_4_22, A1=>nx9348, S0=>nx42609);
   ix9349 : nor02ii port map ( Y=>nx9348, A0=>nx36603, A1=>nx42613);
   ix9343 : xor2 port map ( Y=>nx18386, A0=>nx36622, A1=>nx36779);
   ix9331 : xor2 port map ( Y=>nx18387, A0=>nx36653, A1=>nx42621);
   ix24962 : mux21_ni port map ( Y=>nx24961, A0=>
      booth_booth_integration_output_4_24, A1=>nx9324, S0=>nx42609);
   ix9325 : nor02ii port map ( Y=>nx9324, A0=>nx36639, A1=>nx42613);
   ix9319 : xor2 port map ( Y=>nx18388, A0=>nx36658, A1=>nx36776);
   ix9307 : xor2 port map ( Y=>nx18389, A0=>nx36689, A1=>nx42623);
   ix24942 : mux21_ni port map ( Y=>nx24941, A0=>
      booth_booth_integration_output_4_26, A1=>nx9300, S0=>nx42609);
   ix9301 : nor02ii port map ( Y=>nx9300, A0=>nx36675, A1=>nx42613);
   ix9295 : xor2 port map ( Y=>nx18390, A0=>nx36694, A1=>nx36773);
   ix9283 : xor2 port map ( Y=>nx18391, A0=>nx36725, A1=>nx42625);
   ix24922 : mux21_ni port map ( Y=>nx24921, A0=>booth_output_28_dup_12175, 
      A1=>nx9276, S0=>nx42609);
   ix9277 : nor02ii port map ( Y=>nx9276, A0=>nx36711, A1=>nx42613);
   ix9271 : xor2 port map ( Y=>nx18393, A0=>nx36730, A1=>nx36770);
   ix9259 : xor2 port map ( Y=>nx18395, A0=>nx36746, A1=>nx42627);
   ix36764 : xor2 port map ( Y=>nx36763, A0=>nx36746, A1=>nx9244);
   ix9433 : nor02ii port map ( Y=>nx9432, A0=>nx8896, A1=>nx42613);
   ix36800 : xnor2 port map ( Y=>nx36799, A0=>nx36795, A1=>nx36809);
   ix25122 : mux21_ni port map ( Y=>nx25121, A0=>label_5_output_1, A1=>
      label_5_input_1, S0=>nx43423);
   ix9523 : mux21_ni port map ( Y=>nx9522, A0=>nx9518, A1=>
      label_5_input_state_machine_1, S0=>nx43077);
   ix25112 : mux21_ni port map ( Y=>nx25111, A0=>
      label_5_input_state_machine_1, A1=>data_in(65), S0=>nx42797);
   ix36815 : xnor2 port map ( Y=>nx36814, A0=>nx36792, A1=>nx36824);
   ix25162 : mux21_ni port map ( Y=>nx25161, A0=>label_5_output_3, A1=>
      label_5_input_3, S0=>nx43423);
   ix9587 : mux21_ni port map ( Y=>nx9586, A0=>nx9582, A1=>
      label_5_input_state_machine_3, S0=>nx43079);
   ix25152 : mux21_ni port map ( Y=>nx25151, A0=>
      label_5_input_state_machine_3, A1=>data_in(67), S0=>nx42797);
   ix36826 : xor2 port map ( Y=>nx36825, A0=>nx36499, A1=>label_5_output_4);
   ix36830 : xnor2 port map ( Y=>nx36829, A0=>nx36509, A1=>nx36839);
   ix25202 : mux21_ni port map ( Y=>nx25201, A0=>label_5_output_5, A1=>
      label_5_input_5, S0=>nx43423);
   ix9651 : mux21_ni port map ( Y=>nx9650, A0=>nx9646, A1=>
      label_5_input_state_machine_5, S0=>nx43079);
   ix25192 : mux21_ni port map ( Y=>nx25191, A0=>
      label_5_input_state_machine_5, A1=>data_in(69), S0=>nx42797);
   ix36841 : xor2 port map ( Y=>nx36840, A0=>nx36529, A1=>label_5_output_6);
   ix36845 : xnor2 port map ( Y=>nx36844, A0=>nx36548, A1=>nx36854);
   ix25242 : mux21_ni port map ( Y=>nx25241, A0=>label_5_output_7, A1=>
      label_5_input_7, S0=>nx43423);
   ix9715 : mux21_ni port map ( Y=>nx9714, A0=>nx9710, A1=>
      label_5_input_state_machine_7, S0=>nx43079);
   ix25232 : mux21_ni port map ( Y=>nx25231, A0=>
      label_5_input_state_machine_7, A1=>data_in(71), S0=>nx42797);
   ix36856 : xor2 port map ( Y=>nx36855, A0=>nx36581, A1=>label_5_output_8);
   ix36860 : xnor2 port map ( Y=>nx36859, A0=>nx36586, A1=>nx36869);
   ix25282 : mux21_ni port map ( Y=>nx25281, A0=>label_5_output_9, A1=>
      label_5_input_9, S0=>nx43423);
   ix9779 : mux21_ni port map ( Y=>nx9778, A0=>nx9774, A1=>
      label_5_input_state_machine_9, S0=>nx43079);
   ix25272 : mux21_ni port map ( Y=>nx25271, A0=>
      label_5_input_state_machine_9, A1=>data_in(73), S0=>nx42797);
   ix36871 : xor2 port map ( Y=>nx36870, A0=>nx36617, A1=>label_5_output_10
   );
   ix36875 : xnor2 port map ( Y=>nx36874, A0=>nx36622, A1=>nx36884);
   ix25322 : mux21_ni port map ( Y=>nx25321, A0=>label_5_output_11, A1=>
      label_5_input_11, S0=>nx42811);
   ix9843 : mux21_ni port map ( Y=>nx9842, A0=>nx9838, A1=>
      label_5_input_state_machine_11, S0=>nx43079);
   ix25312 : mux21_ni port map ( Y=>nx25311, A0=>
      label_5_input_state_machine_11, A1=>data_in(75), S0=>nx43373);
   ix36886 : xor2 port map ( Y=>nx36885, A0=>nx36653, A1=>label_5_output_12
   );
   ix36890 : xnor2 port map ( Y=>nx36889, A0=>nx36658, A1=>nx36899);
   ix25362 : mux21_ni port map ( Y=>nx25361, A0=>label_5_output_13, A1=>
      label_5_input_13, S0=>nx42811);
   ix9907 : mux21_ni port map ( Y=>nx9906, A0=>nx9902, A1=>
      label_5_input_state_machine_13, S0=>nx43079);
   ix25352 : mux21_ni port map ( Y=>nx25351, A0=>
      label_5_input_state_machine_13, A1=>data_in(77), S0=>nx43373);
   ix36901 : xor2 port map ( Y=>nx36900, A0=>nx36689, A1=>label_5_output_14
   );
   ix26212 : mux21_ni port map ( Y=>nx26211, A0=>label_6_output_14, A1=>
      label_6_input_14, S0=>nx43425);
   ix11251 : mux21_ni port map ( Y=>nx11250, A0=>nx11246, A1=>
      label_6_input_state_machine_14, S0=>nx43079);
   ix25392 : mux21_ni port map ( Y=>nx25391, A0=>
      label_6_input_state_machine_14, A1=>data_in(94), S0=>nx43373);
   ix26182 : mux21_ni port map ( Y=>nx26181, A0=>label_6_output_12, A1=>
      label_6_input_12, S0=>nx43425);
   ix11193 : mux21_ni port map ( Y=>nx11192, A0=>nx11188, A1=>
      label_6_input_state_machine_12, S0=>nx43081);
   ix26172 : mux21_ni port map ( Y=>nx26171, A0=>
      label_6_input_state_machine_12, A1=>data_in(92), S0=>nx43373);
   ix26142 : mux21_ni port map ( Y=>nx26141, A0=>label_6_output_10, A1=>
      label_6_input_10, S0=>nx43425);
   ix11129 : mux21_ni port map ( Y=>nx11128, A0=>nx11124, A1=>
      label_6_input_state_machine_10, S0=>nx43081);
   ix26132 : mux21_ni port map ( Y=>nx26131, A0=>
      label_6_input_state_machine_10, A1=>data_in(90), S0=>nx43373);
   ix26102 : mux21_ni port map ( Y=>nx26101, A0=>label_6_output_8, A1=>
      label_6_input_8, S0=>nx43425);
   ix11065 : mux21_ni port map ( Y=>nx11064, A0=>nx11060, A1=>
      label_6_input_state_machine_8, S0=>nx43081);
   ix26092 : mux21_ni port map ( Y=>nx26091, A0=>
      label_6_input_state_machine_8, A1=>data_in(88), S0=>nx43373);
   ix26062 : mux21_ni port map ( Y=>nx26061, A0=>label_6_output_6, A1=>
      label_6_input_6, S0=>nx43425);
   ix11001 : mux21_ni port map ( Y=>nx11000, A0=>nx10996, A1=>
      label_6_input_state_machine_6, S0=>nx43081);
   ix26052 : mux21_ni port map ( Y=>nx26051, A0=>
      label_6_input_state_machine_6, A1=>data_in(86), S0=>nx43373);
   ix26022 : mux21_ni port map ( Y=>nx26021, A0=>label_6_output_4, A1=>
      label_6_input_4, S0=>nx42811);
   ix10937 : mux21_ni port map ( Y=>nx10936, A0=>nx10932, A1=>
      label_6_input_state_machine_4, S0=>nx43081);
   ix26012 : mux21_ni port map ( Y=>nx26011, A0=>
      label_6_input_state_machine_4, A1=>data_in(84), S0=>nx43375);
   ix25982 : mux21_ni port map ( Y=>nx25981, A0=>label_6_output_2, A1=>
      label_6_input_2, S0=>nx42811);
   ix10873 : mux21_ni port map ( Y=>nx10872, A0=>nx10868, A1=>
      label_6_input_state_machine_2, S0=>nx43081);
   ix25972 : mux21_ni port map ( Y=>nx25971, A0=>
      label_6_input_state_machine_2, A1=>data_in(82), S0=>nx43375);
   ix25942 : mux21_ni port map ( Y=>nx25941, A0=>label_6_output_0, A1=>
      label_6_input_0, S0=>nx42811);
   ix25932 : mux21_ni port map ( Y=>nx25931, A0=>
      label_6_input_state_machine_0, A1=>data_in(80), S0=>nx43375);
   ix25922 : mux21_ni port map ( Y=>nx25921, A0=>
      booth_booth_integration_output_5_12, A1=>nx10792, S0=>nx43269);
   ix10793 : mux21_ni port map ( Y=>nx10792, A0=>nx41809, A1=>
      booth_booth_integration_output_5_13, S0=>nx43277);
   ix25912 : mux21_ni port map ( Y=>nx25911, A0=>
      booth_booth_integration_output_5_13, A1=>nx10780, S0=>nx43269);
   ix10781 : mux21_ni port map ( Y=>nx10780, A0=>nx41805, A1=>
      booth_booth_integration_output_5_14, S0=>nx43277);
   ix25902 : mux21_ni port map ( Y=>nx25901, A0=>
      booth_booth_integration_output_5_14, A1=>nx10768, S0=>nx43269);
   ix10769 : mux21_ni port map ( Y=>nx10768, A0=>nx41801, A1=>
      booth_booth_integration_output_5_15, S0=>nx43277);
   ix25892 : mux21 port map ( Y=>nx25891, A0=>nx37428, A1=>nx37009, S0=>
      nx43269);
   ix25422 : mux21_ni port map ( Y=>nx25421, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_0, A1=>nx42015, S0=>nx42949
   );
   ix25408 : and02 port map ( Y=>nx25407, A0=>nx43487, A1=>
      booth_booth_integrtaion_5_shift_Reg_count_0);
   ix25602 : mux21_ni port map ( Y=>nx25601, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_9, A1=>nx42001, S0=>nx42949
   );
   ix25592 : mux21_ni port map ( Y=>nx25591, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_9, A1=>output_8_dup_12828, 
      S0=>nx43269);
   ix25582 : mux21_ni port map ( Y=>nx25581, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_8, A1=>output_8_dup_12828, 
      S0=>nx42949);
   ix25572 : mux21_ni port map ( Y=>nx25571, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_8, A1=>output_7_dup_12829, 
      S0=>nx43269);
   ix25562 : mux21_ni port map ( Y=>nx25561, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_7, A1=>output_7_dup_12829, 
      S0=>nx42949);
   ix25552 : mux21_ni port map ( Y=>nx25551, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_7, A1=>output_6_dup_12830, 
      S0=>nx43271);
   ix25542 : mux21_ni port map ( Y=>nx25541, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_6, A1=>output_6_dup_12830, 
      S0=>nx42949);
   ix25532 : mux21_ni port map ( Y=>nx25531, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_6, A1=>output_5_dup_12831, 
      S0=>nx43271);
   ix25522 : mux21_ni port map ( Y=>nx25521, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_5, A1=>output_5_dup_12831, 
      S0=>nx42949);
   ix25512 : mux21_ni port map ( Y=>nx25511, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_5, A1=>output_4_dup_12832, 
      S0=>nx43271);
   ix25502 : mux21_ni port map ( Y=>nx25501, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_4, A1=>output_4_dup_12832, 
      S0=>nx42951);
   ix25492 : mux21_ni port map ( Y=>nx25491, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_4, A1=>output_3_dup_12833, 
      S0=>nx43271);
   ix25482 : mux21_ni port map ( Y=>nx25481, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_3, A1=>output_3_dup_12833, 
      S0=>nx42951);
   ix25472 : mux21_ni port map ( Y=>nx25471, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_3, A1=>output_2_dup_12834, 
      S0=>nx43271);
   ix25462 : mux21_ni port map ( Y=>nx25461, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_2, A1=>output_2_dup_12834, 
      S0=>nx42951);
   ix25452 : mux21_ni port map ( Y=>nx25451, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_2, A1=>output_1_dup_12835, 
      S0=>nx43271);
   ix25442 : mux21_ni port map ( Y=>nx25441, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_1, A1=>output_1_dup_12835, 
      S0=>nx42951);
   ix25432 : mux21_ni port map ( Y=>nx25431, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_1, A1=>nx42015, S0=>nx43271
   );
   ix10209 : nand02 port map ( Y=>nx37155, A0=>nx37082, A1=>
      booth_output_0_dup_12206);
   ix37085 : or03 port map ( Y=>nx37084, A0=>nx37133, A1=>
      booth_booth_integrtaion_5_shift_reg_output_0, A2=>nx43487);
   ix25722 : mux21_ni port map ( Y=>nx25721, A0=>booth_output_0_dup_12206, 
      A1=>nx10188, S0=>nx43273);
   ix10189 : mux21_ni port map ( Y=>nx10188, A0=>nx41783, A1=>
      booth_output_1_dup_12205, S0=>nx43279);
   ix25712 : mux21_ni port map ( Y=>nx25711, A0=>booth_output_1_dup_12205, 
      A1=>nx10176, S0=>nx43273);
   ix10177 : mux21_ni port map ( Y=>nx10176, A0=>nx41779, A1=>
      booth_output_2_dup_12204, S0=>nx43279);
   ix25702 : mux21_ni port map ( Y=>nx25701, A0=>booth_output_2_dup_12204, 
      A1=>nx10164, S0=>nx43273);
   ix10165 : mux21_ni port map ( Y=>nx10164, A0=>nx41775, A1=>
      booth_output_3_dup_12203, S0=>nx43279);
   ix25692 : mux21_ni port map ( Y=>nx25691, A0=>booth_output_3_dup_12203, 
      A1=>nx10152, S0=>nx43273);
   ix10153 : mux21_ni port map ( Y=>nx10152, A0=>nx41771, A1=>
      booth_output_4_dup_12202, S0=>nx43279);
   ix25682 : mux21_ni port map ( Y=>nx25681, A0=>booth_output_4_dup_12202, 
      A1=>nx10140, S0=>nx43273);
   ix10141 : mux21_ni port map ( Y=>nx10140, A0=>nx41767, A1=>
      booth_output_5_dup_12201, S0=>nx43279);
   ix25672 : mux21_ni port map ( Y=>nx25671, A0=>booth_output_5_dup_12201, 
      A1=>nx10128, S0=>nx43273);
   ix10129 : mux21_ni port map ( Y=>nx10128, A0=>nx41763, A1=>
      booth_output_6_dup_12200, S0=>nx43279);
   ix25662 : mux21_ni port map ( Y=>nx25661, A0=>booth_output_6_dup_12200, 
      A1=>nx10116, S0=>nx43273);
   ix10117 : mux21_ni port map ( Y=>nx10116, A0=>nx41759, A1=>
      booth_output_7_dup_12199, S0=>nx43279);
   ix25652 : mux21_ni port map ( Y=>nx25651, A0=>booth_output_7_dup_12199, 
      A1=>nx10104, S0=>nx43275);
   ix10105 : mux21_ni port map ( Y=>nx10104, A0=>nx41755, A1=>
      booth_output_8_dup_12198, S0=>nx43281);
   ix25642 : mux21_ni port map ( Y=>nx25641, A0=>booth_output_8_dup_12198, 
      A1=>nx10092, S0=>nx43275);
   ix10093 : mux21_ni port map ( Y=>nx10092, A0=>nx41751, A1=>
      booth_output_9_dup_12197, S0=>nx43281);
   ix25632 : mux21_ni port map ( Y=>nx25631, A0=>booth_output_9_dup_12197, 
      A1=>nx10080, S0=>nx43275);
   ix10081 : mux21_ni port map ( Y=>nx10080, A0=>nx41747, A1=>
      booth_output_10_dup_12196, S0=>nx43281);
   ix25622 : mux21_ni port map ( Y=>nx25621, A0=>booth_output_10_dup_12196, 
      A1=>nx10068, S0=>nx43275);
   ix10069 : mux21_ni port map ( Y=>nx10068, A0=>nx41743, A1=>
      booth_output_11_dup_12195, S0=>nx43281);
   ix25612 : mux21_ni port map ( Y=>nx25611, A0=>booth_output_11_dup_12195, 
      A1=>nx10056, S0=>nx43275);
   ix10057 : mux21_ni port map ( Y=>nx10056, A0=>nx41731, A1=>
      booth_booth_integration_output_5_12, S0=>nx43281);
   ix25882 : mux21_ni port map ( Y=>nx25881, A0=>
      booth_booth_integration_output_5_16, A1=>nx10738, S0=>nx43275);
   ix10739 : nor02ii port map ( Y=>nx10738, A0=>nx37139, A1=>nx43281);
   ix10215 : nor02ii port map ( Y=>nx10214, A0=>nx37077, A1=>
      booth_booth_integration_output_5_16);
   ix10733 : xor2 port map ( Y=>nx18421, A0=>nx37145, A1=>nx37421);
   ix37161 : or02 port map ( Y=>nx37160, A0=>nx37082, A1=>
      booth_output_0_dup_12206);
   ix10721 : xor2 port map ( Y=>nx18422, A0=>nx37165, A1=>nx42663);
   ix37181 : xor2 port map ( Y=>nx37180, A0=>nx37184, A1=>nx10286);
   ix37193 : nor02ii port map ( Y=>nx37192, A0=>nx10252, A1=>data_in(83));
   ix10697 : xor2 port map ( Y=>nx18424, A0=>nx37217, A1=>nx42665);
   ix25842 : mux21_ni port map ( Y=>nx25841, A0=>
      booth_booth_integration_output_5_20, A1=>nx10690, S0=>nx43275);
   ix10691 : nor02ii port map ( Y=>nx10690, A0=>nx37203, A1=>nx43281);
   ix10685 : xor2 port map ( Y=>nx18425, A0=>nx37222, A1=>nx37418);
   ix10673 : xor2 port map ( Y=>nx18426, A0=>nx37253, A1=>nx42667);
   ix25822 : mux21_ni port map ( Y=>nx25821, A0=>
      booth_booth_integration_output_5_22, A1=>nx10666, S0=>nx42657);
   ix10667 : nor02ii port map ( Y=>nx10666, A0=>nx37239, A1=>nx42661);
   ix10661 : xor2 port map ( Y=>nx18427, A0=>nx37258, A1=>nx37415);
   ix10649 : xor2 port map ( Y=>nx18429, A0=>nx37289, A1=>nx42669);
   ix25802 : mux21_ni port map ( Y=>nx25801, A0=>
      booth_booth_integration_output_5_24, A1=>nx10642, S0=>nx42657);
   ix10643 : nor02ii port map ( Y=>nx10642, A0=>nx37275, A1=>nx42661);
   ix10637 : xor2 port map ( Y=>nx18431, A0=>nx37294, A1=>nx37412);
   ix10625 : xor2 port map ( Y=>nx18433, A0=>nx37325, A1=>nx42671);
   ix25782 : mux21_ni port map ( Y=>nx25781, A0=>
      booth_booth_integration_output_5_26, A1=>nx10618, S0=>nx42657);
   ix10619 : nor02ii port map ( Y=>nx10618, A0=>nx37311, A1=>nx42661);
   ix10613 : xor2 port map ( Y=>nx18435, A0=>nx37330, A1=>nx37409);
   ix10601 : xor2 port map ( Y=>nx18437, A0=>nx37361, A1=>nx42673);
   ix25762 : mux21_ni port map ( Y=>nx25761, A0=>booth_output_28_dup_12194, 
      A1=>nx10594, S0=>nx42657);
   ix10595 : nor02ii port map ( Y=>nx10594, A0=>nx37347, A1=>nx42661);
   ix10589 : xor2 port map ( Y=>nx18439, A0=>nx37366, A1=>nx37406);
   ix10577 : xor2 port map ( Y=>nx18440, A0=>nx37382, A1=>nx42675);
   ix37400 : xor2 port map ( Y=>nx37399, A0=>nx37382, A1=>nx10562);
   ix10751 : nor02ii port map ( Y=>nx10750, A0=>nx10214, A1=>nx42661);
   ix37436 : xnor2 port map ( Y=>nx37435, A0=>nx37431, A1=>nx37445);
   ix25962 : mux21_ni port map ( Y=>nx25961, A0=>label_6_output_1, A1=>
      label_6_input_1, S0=>nx42811);
   ix10841 : mux21_ni port map ( Y=>nx10840, A0=>nx10836, A1=>
      label_6_input_state_machine_1, S0=>nx43081);
   ix25952 : mux21_ni port map ( Y=>nx25951, A0=>
      label_6_input_state_machine_1, A1=>data_in(81), S0=>nx43375);
   ix37451 : xnor2 port map ( Y=>nx37450, A0=>nx37428, A1=>nx37460);
   ix26002 : mux21_ni port map ( Y=>nx26001, A0=>label_6_output_3, A1=>
      label_6_input_3, S0=>nx42811);
   ix10905 : mux21_ni port map ( Y=>nx10904, A0=>nx10900, A1=>
      label_6_input_state_machine_3, S0=>nx43083);
   ix25992 : mux21_ni port map ( Y=>nx25991, A0=>
      label_6_input_state_machine_3, A1=>data_in(83), S0=>nx43375);
   ix37462 : xor2 port map ( Y=>nx37461, A0=>nx37135, A1=>label_6_output_4);
   ix37466 : xnor2 port map ( Y=>nx37465, A0=>nx37145, A1=>nx37475);
   ix26042 : mux21_ni port map ( Y=>nx26041, A0=>label_6_output_5, A1=>
      label_6_input_5, S0=>nx43425);
   ix10969 : mux21_ni port map ( Y=>nx10968, A0=>nx10964, A1=>
      label_6_input_state_machine_5, S0=>nx43083);
   ix26032 : mux21_ni port map ( Y=>nx26031, A0=>
      label_6_input_state_machine_5, A1=>data_in(85), S0=>nx43375);
   ix37477 : xor2 port map ( Y=>nx37476, A0=>nx37165, A1=>label_6_output_6);
   ix37481 : xnor2 port map ( Y=>nx37480, A0=>nx37184, A1=>nx37490);
   ix26082 : mux21_ni port map ( Y=>nx26081, A0=>label_6_output_7, A1=>
      label_6_input_7, S0=>nx43425);
   ix11033 : mux21_ni port map ( Y=>nx11032, A0=>nx11028, A1=>
      label_6_input_state_machine_7, S0=>nx43083);
   ix26072 : mux21_ni port map ( Y=>nx26071, A0=>
      label_6_input_state_machine_7, A1=>data_in(87), S0=>nx43375);
   ix37492 : xor2 port map ( Y=>nx37491, A0=>nx37217, A1=>label_6_output_8);
   ix37496 : xnor2 port map ( Y=>nx37495, A0=>nx37222, A1=>nx37505);
   ix26122 : mux21_ni port map ( Y=>nx26121, A0=>label_6_output_9, A1=>
      label_6_input_9, S0=>nx43427);
   ix11097 : mux21_ni port map ( Y=>nx11096, A0=>nx11092, A1=>
      label_6_input_state_machine_9, S0=>nx43083);
   ix26112 : mux21_ni port map ( Y=>nx26111, A0=>
      label_6_input_state_machine_9, A1=>data_in(89), S0=>nx43377);
   ix37507 : xor2 port map ( Y=>nx37506, A0=>nx37253, A1=>label_6_output_10
   );
   ix37511 : xnor2 port map ( Y=>nx37510, A0=>nx37258, A1=>nx37520);
   ix26162 : mux21_ni port map ( Y=>nx26161, A0=>label_6_output_11, A1=>
      label_6_input_11, S0=>nx43427);
   ix11161 : mux21_ni port map ( Y=>nx11160, A0=>nx11156, A1=>
      label_6_input_state_machine_11, S0=>nx43083);
   ix26152 : mux21_ni port map ( Y=>nx26151, A0=>
      label_6_input_state_machine_11, A1=>data_in(91), S0=>nx43377);
   ix37522 : xor2 port map ( Y=>nx37521, A0=>nx37289, A1=>label_6_output_12
   );
   ix37526 : xnor2 port map ( Y=>nx37525, A0=>nx37294, A1=>nx37535);
   ix26202 : mux21_ni port map ( Y=>nx26201, A0=>label_6_output_13, A1=>
      label_6_input_13, S0=>nx43427);
   ix11225 : mux21_ni port map ( Y=>nx11224, A0=>nx11220, A1=>
      label_6_input_state_machine_13, S0=>nx43083);
   ix26192 : mux21_ni port map ( Y=>nx26191, A0=>
      label_6_input_state_machine_13, A1=>data_in(93), S0=>nx43377);
   ix37537 : xor2 port map ( Y=>nx37536, A0=>nx37325, A1=>label_6_output_14
   );
   ix11273 : xnor2 port map ( Y=>nx11272, A0=>nx36907, A1=>nx36271);
   ix37545 : xnor2 port map ( Y=>nx37544, A0=>nx37548, A1=>
      max_calc_comparator_third_inp1_13);
   ix37551 : or03 port map ( Y=>nx37550, A0=>nx37535, A1=>nx43341, A2=>
      nx43211);
   ix37556 : or03 port map ( Y=>nx37555, A0=>nx36899, A1=>nx43341, A2=>
      nx43211);
   ix11317 : xnor2 port map ( Y=>nx11316, A0=>nx37559, A1=>nx37566);
   ix37573 : xnor2 port map ( Y=>nx37572, A0=>nx37576, A1=>
      max_calc_comparator_third_inp1_11);
   ix37579 : or03 port map ( Y=>nx37578, A0=>nx37520, A1=>nx43343, A2=>
      nx43211);
   ix37584 : or03 port map ( Y=>nx37583, A0=>nx36884, A1=>nx43343, A2=>
      nx43211);
   ix11361 : xnor2 port map ( Y=>nx11360, A0=>nx37587, A1=>nx37594);
   ix37601 : xnor2 port map ( Y=>nx37600, A0=>nx37604, A1=>
      max_calc_comparator_third_inp1_9);
   ix37607 : or03 port map ( Y=>nx37606, A0=>nx37505, A1=>nx43343, A2=>
      nx43211);
   ix37612 : or03 port map ( Y=>nx37611, A0=>nx36869, A1=>nx43343, A2=>
      nx43211);
   ix11405 : xnor2 port map ( Y=>nx11404, A0=>nx37615, A1=>nx37622);
   ix37629 : xnor2 port map ( Y=>nx37628, A0=>nx37632, A1=>
      max_calc_comparator_third_inp1_7);
   ix37635 : or03 port map ( Y=>nx37634, A0=>nx37490, A1=>nx43343, A2=>
      nx43211);
   ix37640 : or03 port map ( Y=>nx37639, A0=>nx36854, A1=>nx43343, A2=>
      nx42543);
   ix11449 : xnor2 port map ( Y=>nx11448, A0=>nx37643, A1=>nx37650);
   ix37657 : xnor2 port map ( Y=>nx37656, A0=>nx37660, A1=>
      max_calc_comparator_third_inp1_5);
   ix37663 : or03 port map ( Y=>nx37662, A0=>nx37475, A1=>nx43343, A2=>
      nx42543);
   ix37668 : or03 port map ( Y=>nx37667, A0=>nx36839, A1=>nx43345, A2=>
      nx42543);
   ix11493 : xnor2 port map ( Y=>nx11492, A0=>nx37671, A1=>nx37678);
   ix37685 : xnor2 port map ( Y=>nx37684, A0=>nx37688, A1=>
      max_calc_comparator_third_inp1_3);
   ix37691 : or03 port map ( Y=>nx37690, A0=>nx37460, A1=>nx43345, A2=>
      nx42543);
   ix37696 : or03 port map ( Y=>nx37695, A0=>nx36824, A1=>nx43345, A2=>
      nx42543);
   ix11537 : xnor2 port map ( Y=>nx11536, A0=>nx37699, A1=>nx37706);
   ix37717 : or03 port map ( Y=>nx37716, A0=>nx37445, A1=>nx43345, A2=>
      nx42543);
   ix37722 : or03 port map ( Y=>nx37721, A0=>nx36809, A1=>nx43345, A2=>
      nx43215);
   ix11559 : xnor2 port map ( Y=>nx11558, A0=>nx37714, A1=>nx37718);
   ix11785 : xnor2 port map ( Y=>nx11784, A0=>nx37740, A1=>nx37760);
   ix37743 : or03 port map ( Y=>nx37742, A0=>nx37756, A1=>nx43345, A2=>
      nx43215);
   ix26522 : mux21_ni port map ( Y=>nx26521, A0=>label_6_output_15, A1=>
      label_6_input_15, S0=>nx43427);
   ix11721 : mux21_ni port map ( Y=>nx11720, A0=>nx11716, A1=>
      label_6_input_state_machine_15, S0=>nx43083);
   ix26512 : mux21_ni port map ( Y=>nx26511, A0=>
      label_6_input_state_machine_15, A1=>data_in(95), S0=>nx43377);
   ix11715 : xnor2 port map ( Y=>nx11714, A0=>nx37330, A1=>label_6_output_15
   );
   ix37763 : or03 port map ( Y=>nx37762, A0=>nx37776, A1=>nx43345, A2=>
      nx43215);
   ix26552 : mux21_ni port map ( Y=>nx26551, A0=>label_5_output_15, A1=>
      label_5_input_15, S0=>nx43427);
   ix11763 : mux21_ni port map ( Y=>nx11762, A0=>nx11758, A1=>
      label_5_input_state_machine_15, S0=>nx42291);
   ix26542 : mux21_ni port map ( Y=>nx26541, A0=>
      label_5_input_state_machine_15, A1=>data_in(79), S0=>nx43377);
   ix11757 : xnor2 port map ( Y=>nx11756, A0=>nx36694, A1=>label_5_output_15
   );
   ix37779 : nor02_2x port map ( Y=>nx42677, A0=>nx43203, A1=>nx43285);
   ix37781 : nor03_2x port map ( Y=>nx42689, A0=>nx43203, A1=>nx43139, A2=>
      nx42843);
   ix16299 : mux21_ni port map ( Y=>nx16298, A0=>max_calc_ans4_14, A1=>
      label_4_output_14, S0=>nx43139);
   ix27412 : mux21_ni port map ( Y=>nx27411, A0=>label_4_output_14, A1=>
      label_4_input_14, S0=>nx43427);
   ix13115 : mux21_ni port map ( Y=>nx13114, A0=>nx13110, A1=>
      label_4_input_state_machine_14, S0=>nx43085);
   ix26592 : mux21_ni port map ( Y=>nx26591, A0=>
      label_4_input_state_machine_14, A1=>data_in(62), S0=>nx43377);
   ix27382 : mux21_ni port map ( Y=>nx27381, A0=>label_4_output_12, A1=>
      label_4_input_12, S0=>nx43427);
   ix13057 : mux21_ni port map ( Y=>nx13056, A0=>nx13052, A1=>
      label_4_input_state_machine_12, S0=>nx43085);
   ix27372 : mux21_ni port map ( Y=>nx27371, A0=>
      label_4_input_state_machine_12, A1=>data_in(60), S0=>nx43377);
   ix27342 : mux21_ni port map ( Y=>nx27341, A0=>label_4_output_10, A1=>
      label_4_input_10, S0=>nx43429);
   ix12993 : mux21_ni port map ( Y=>nx12992, A0=>nx12988, A1=>
      label_4_input_state_machine_10, S0=>nx43085);
   ix27332 : mux21_ni port map ( Y=>nx27331, A0=>
      label_4_input_state_machine_10, A1=>data_in(58), S0=>nx43379);
   ix27302 : mux21_ni port map ( Y=>nx27301, A0=>label_4_output_8, A1=>
      label_4_input_8, S0=>nx43429);
   ix12929 : mux21_ni port map ( Y=>nx12928, A0=>nx12924, A1=>
      label_4_input_state_machine_8, S0=>nx43085);
   ix27292 : mux21_ni port map ( Y=>nx27291, A0=>
      label_4_input_state_machine_8, A1=>data_in(56), S0=>nx43379);
   ix27262 : mux21_ni port map ( Y=>nx27261, A0=>label_4_output_6, A1=>
      label_4_input_6, S0=>nx43429);
   ix12865 : mux21_ni port map ( Y=>nx12864, A0=>nx12860, A1=>
      label_4_input_state_machine_6, S0=>nx42291);
   ix27252 : mux21_ni port map ( Y=>nx27251, A0=>
      label_4_input_state_machine_6, A1=>data_in(54), S0=>nx43379);
   ix27222 : mux21_ni port map ( Y=>nx27221, A0=>label_4_output_4, A1=>
      label_4_input_4, S0=>nx43429);
   ix12801 : mux21_ni port map ( Y=>nx12800, A0=>nx12796, A1=>
      label_4_input_state_machine_4, S0=>nx42291);
   ix27212 : mux21_ni port map ( Y=>nx27211, A0=>
      label_4_input_state_machine_4, A1=>data_in(52), S0=>nx43379);
   ix27182 : mux21_ni port map ( Y=>nx27181, A0=>label_4_output_2, A1=>
      label_4_input_2, S0=>nx43429);
   ix12737 : mux21_ni port map ( Y=>nx12736, A0=>nx12732, A1=>
      label_4_input_state_machine_2, S0=>nx42291);
   ix27172 : mux21_ni port map ( Y=>nx27171, A0=>
      label_4_input_state_machine_2, A1=>data_in(50), S0=>nx43379);
   ix27142 : mux21_ni port map ( Y=>nx27141, A0=>label_4_output_0, A1=>
      label_4_input_0, S0=>nx43429);
   ix27132 : mux21_ni port map ( Y=>nx27131, A0=>
      label_4_input_state_machine_0, A1=>data_in(48), S0=>nx43379);
   ix27122 : mux21_ni port map ( Y=>nx27121, A0=>
      booth_booth_integration_output_3_12, A1=>nx12656, S0=>nx43291);
   ix12657 : mux21_ni port map ( Y=>nx12656, A0=>nx41809, A1=>
      booth_booth_integration_output_3_13, S0=>nx43299);
   ix27112 : mux21_ni port map ( Y=>nx27111, A0=>
      booth_booth_integration_output_3_13, A1=>nx12644, S0=>nx43291);
   ix12645 : mux21_ni port map ( Y=>nx12644, A0=>nx41805, A1=>
      booth_booth_integration_output_3_14, S0=>nx43299);
   ix27102 : mux21_ni port map ( Y=>nx27101, A0=>
      booth_booth_integration_output_3_14, A1=>nx12632, S0=>nx43291);
   ix12633 : mux21_ni port map ( Y=>nx12632, A0=>nx41801, A1=>
      booth_booth_integration_output_3_15, S0=>nx43299);
   ix27092 : mux21 port map ( Y=>nx27091, A0=>nx38307, A1=>nx37888, S0=>
      nx43291);
   ix26622 : mux21_ni port map ( Y=>nx26621, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_0, A1=>nx42055, S0=>nx42953
   );
   ix26608 : and02 port map ( Y=>nx26607, A0=>nx43491, A1=>
      booth_booth_integrtaion_3_shift_Reg_count_0);
   ix26802 : mux21_ni port map ( Y=>nx26801, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_9, A1=>nx42041, S0=>nx42953
   );
   ix26792 : mux21_ni port map ( Y=>nx26791, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_9, A1=>output_8_dup_12772, 
      S0=>nx43291);
   ix26782 : mux21_ni port map ( Y=>nx26781, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_8, A1=>output_8_dup_12772, 
      S0=>nx42953);
   ix26772 : mux21_ni port map ( Y=>nx26771, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_8, A1=>output_7_dup_12773, 
      S0=>nx43291);
   ix26762 : mux21_ni port map ( Y=>nx26761, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_7, A1=>output_7_dup_12773, 
      S0=>nx42953);
   ix26752 : mux21_ni port map ( Y=>nx26751, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_7, A1=>output_6_dup_12774, 
      S0=>nx43293);
   ix26742 : mux21_ni port map ( Y=>nx26741, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_6, A1=>output_6_dup_12774, 
      S0=>nx42953);
   ix26732 : mux21_ni port map ( Y=>nx26731, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_6, A1=>output_5_dup_12775, 
      S0=>nx43293);
   ix26722 : mux21_ni port map ( Y=>nx26721, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_5, A1=>output_5_dup_12775, 
      S0=>nx42953);
   ix26712 : mux21_ni port map ( Y=>nx26711, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_5, A1=>output_4_dup_12776, 
      S0=>nx43293);
   ix26702 : mux21_ni port map ( Y=>nx26701, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_4, A1=>output_4_dup_12776, 
      S0=>nx42955);
   ix26692 : mux21_ni port map ( Y=>nx26691, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_4, A1=>output_3_dup_12777, 
      S0=>nx43293);
   ix26682 : mux21_ni port map ( Y=>nx26681, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_3, A1=>output_3_dup_12777, 
      S0=>nx42955);
   ix26672 : mux21_ni port map ( Y=>nx26671, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_3, A1=>output_2_dup_12778, 
      S0=>nx43293);
   ix26662 : mux21_ni port map ( Y=>nx26661, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_2, A1=>output_2_dup_12778, 
      S0=>nx42955);
   ix26652 : mux21_ni port map ( Y=>nx26651, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_2, A1=>output_1_dup_12779, 
      S0=>nx43293);
   ix26642 : mux21_ni port map ( Y=>nx26641, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_1, A1=>output_1_dup_12779, 
      S0=>nx42955);
   ix26632 : mux21_ni port map ( Y=>nx26631, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_1, A1=>nx42055, S0=>nx43293
   );
   ix12073 : nand02 port map ( Y=>nx38034, A0=>nx37961, A1=>
      booth_output_0_dup_12168);
   ix37964 : or03 port map ( Y=>nx37963, A0=>nx38012, A1=>
      booth_booth_integrtaion_3_shift_reg_output_0, A2=>nx43491);
   ix26922 : mux21_ni port map ( Y=>nx26921, A0=>booth_output_0_dup_12168, 
      A1=>nx12052, S0=>nx43295);
   ix12053 : mux21_ni port map ( Y=>nx12052, A0=>nx41783, A1=>
      booth_output_1_dup_12167, S0=>nx43301);
   ix26912 : mux21_ni port map ( Y=>nx26911, A0=>booth_output_1_dup_12167, 
      A1=>nx12040, S0=>nx43295);
   ix12041 : mux21_ni port map ( Y=>nx12040, A0=>nx41779, A1=>
      booth_output_2_dup_12166, S0=>nx43301);
   ix26902 : mux21_ni port map ( Y=>nx26901, A0=>booth_output_2_dup_12166, 
      A1=>nx12028, S0=>nx43295);
   ix12029 : mux21_ni port map ( Y=>nx12028, A0=>nx41775, A1=>
      booth_output_3_dup_12165, S0=>nx43301);
   ix26892 : mux21_ni port map ( Y=>nx26891, A0=>booth_output_3_dup_12165, 
      A1=>nx12016, S0=>nx43295);
   ix12017 : mux21_ni port map ( Y=>nx12016, A0=>nx41771, A1=>
      booth_output_4_dup_12164, S0=>nx43301);
   ix26882 : mux21_ni port map ( Y=>nx26881, A0=>booth_output_4_dup_12164, 
      A1=>nx12004, S0=>nx43295);
   ix12005 : mux21_ni port map ( Y=>nx12004, A0=>nx41767, A1=>
      booth_output_5_dup_12163, S0=>nx43301);
   ix26872 : mux21_ni port map ( Y=>nx26871, A0=>booth_output_5_dup_12163, 
      A1=>nx11992, S0=>nx43295);
   ix11993 : mux21_ni port map ( Y=>nx11992, A0=>nx41763, A1=>
      booth_output_6_dup_12162, S0=>nx43301);
   ix26862 : mux21_ni port map ( Y=>nx26861, A0=>booth_output_6_dup_12162, 
      A1=>nx11980, S0=>nx43295);
   ix11981 : mux21_ni port map ( Y=>nx11980, A0=>nx41759, A1=>
      booth_output_7_dup_12161, S0=>nx43301);
   ix26852 : mux21_ni port map ( Y=>nx26851, A0=>booth_output_7_dup_12161, 
      A1=>nx11968, S0=>nx43297);
   ix11969 : mux21_ni port map ( Y=>nx11968, A0=>nx41755, A1=>
      booth_output_8_dup_12160, S0=>nx43303);
   ix26842 : mux21_ni port map ( Y=>nx26841, A0=>booth_output_8_dup_12160, 
      A1=>nx11956, S0=>nx43297);
   ix11957 : mux21_ni port map ( Y=>nx11956, A0=>nx41751, A1=>
      booth_output_9_dup_12159, S0=>nx43303);
   ix26832 : mux21_ni port map ( Y=>nx26831, A0=>booth_output_9_dup_12159, 
      A1=>nx11944, S0=>nx43297);
   ix11945 : mux21_ni port map ( Y=>nx11944, A0=>nx41747, A1=>
      booth_output_10_dup_12158, S0=>nx43303);
   ix26822 : mux21_ni port map ( Y=>nx26821, A0=>booth_output_10_dup_12158, 
      A1=>nx11932, S0=>nx43297);
   ix11933 : mux21_ni port map ( Y=>nx11932, A0=>nx41743, A1=>
      booth_output_11_dup_12157, S0=>nx43303);
   ix26812 : mux21_ni port map ( Y=>nx26811, A0=>booth_output_11_dup_12157, 
      A1=>nx11920, S0=>nx43297);
   ix11921 : mux21_ni port map ( Y=>nx11920, A0=>nx41731, A1=>
      booth_booth_integration_output_3_12, S0=>nx43303);
   ix27082 : mux21_ni port map ( Y=>nx27081, A0=>
      booth_booth_integration_output_3_16, A1=>nx12602, S0=>nx43297);
   ix12603 : nor02ii port map ( Y=>nx12602, A0=>nx38018, A1=>nx43303);
   ix12079 : nor02ii port map ( Y=>nx12078, A0=>nx37956, A1=>
      booth_booth_integration_output_3_16);
   ix12597 : xor2 port map ( Y=>nx18461, A0=>nx38024, A1=>nx38300);
   ix38040 : or02 port map ( Y=>nx38039, A0=>nx37961, A1=>
      booth_output_0_dup_12168);
   ix12585 : xor2 port map ( Y=>nx18463, A0=>nx38044, A1=>nx42709);
   ix38060 : xor2 port map ( Y=>nx38059, A0=>nx38063, A1=>nx12150);
   ix38072 : nor02ii port map ( Y=>nx38071, A0=>nx12116, A1=>data_in(51));
   ix12561 : xor2 port map ( Y=>nx18467, A0=>nx38096, A1=>nx42711);
   ix27042 : mux21_ni port map ( Y=>nx27041, A0=>
      booth_booth_integration_output_3_20, A1=>nx12554, S0=>nx43297);
   ix12555 : nor02ii port map ( Y=>nx12554, A0=>nx38082, A1=>nx43303);
   ix12549 : xor2 port map ( Y=>nx18469, A0=>nx38101, A1=>nx38297);
   ix12537 : xor2 port map ( Y=>nx18471, A0=>nx38132, A1=>nx42713);
   ix27022 : mux21_ni port map ( Y=>nx27021, A0=>
      booth_booth_integration_output_3_22, A1=>nx12530, S0=>nx42703);
   ix12531 : nor02ii port map ( Y=>nx12530, A0=>nx38118, A1=>nx42707);
   ix12525 : xor2 port map ( Y=>nx18472, A0=>nx38137, A1=>nx38294);
   ix12513 : xor2 port map ( Y=>nx18473, A0=>nx38168, A1=>nx42715);
   ix27002 : mux21_ni port map ( Y=>nx27001, A0=>
      booth_booth_integration_output_3_24, A1=>nx12506, S0=>nx42703);
   ix12507 : nor02ii port map ( Y=>nx12506, A0=>nx38154, A1=>nx42707);
   ix12501 : xor2 port map ( Y=>nx18474, A0=>nx38173, A1=>nx38291);
   ix12489 : xor2 port map ( Y=>nx18475, A0=>nx38204, A1=>nx42717);
   ix26982 : mux21_ni port map ( Y=>nx26981, A0=>
      booth_booth_integration_output_3_26, A1=>nx12482, S0=>nx42703);
   ix12483 : nor02ii port map ( Y=>nx12482, A0=>nx38190, A1=>nx42707);
   ix12477 : xor2 port map ( Y=>nx18476, A0=>nx38209, A1=>nx38288);
   ix12465 : xor2 port map ( Y=>nx18477, A0=>nx38240, A1=>nx42719);
   ix26962 : mux21_ni port map ( Y=>nx26961, A0=>booth_output_28_dup_12156, 
      A1=>nx12458, S0=>nx42703);
   ix12459 : nor02ii port map ( Y=>nx12458, A0=>nx38226, A1=>nx42707);
   ix12453 : xor2 port map ( Y=>nx18479, A0=>nx38245, A1=>nx38285);
   ix12441 : xor2 port map ( Y=>nx18481, A0=>nx38261, A1=>nx42721);
   ix38279 : xor2 port map ( Y=>nx38278, A0=>nx38261, A1=>nx12426);
   ix12615 : nor02ii port map ( Y=>nx12614, A0=>nx12078, A1=>nx42707);
   ix38315 : xnor2 port map ( Y=>nx38314, A0=>nx38310, A1=>nx38324);
   ix27162 : mux21_ni port map ( Y=>nx27161, A0=>label_4_output_1, A1=>
      label_4_input_1, S0=>nx43429);
   ix12705 : mux21_ni port map ( Y=>nx12704, A0=>nx12700, A1=>
      label_4_input_state_machine_1, S0=>nx42291);
   ix27152 : mux21_ni port map ( Y=>nx27151, A0=>
      label_4_input_state_machine_1, A1=>data_in(49), S0=>nx43379);
   ix38330 : xnor2 port map ( Y=>nx38329, A0=>nx38307, A1=>nx38339);
   ix27202 : mux21_ni port map ( Y=>nx27201, A0=>label_4_output_3, A1=>
      label_4_input_3, S0=>nx43431);
   ix12769 : mux21_ni port map ( Y=>nx12768, A0=>nx12764, A1=>
      label_4_input_state_machine_3, S0=>nx42291);
   ix27192 : mux21_ni port map ( Y=>nx27191, A0=>
      label_4_input_state_machine_3, A1=>data_in(51), S0=>nx43381);
   ix38341 : xor2 port map ( Y=>nx38340, A0=>nx38014, A1=>label_4_output_4);
   ix38345 : xnor2 port map ( Y=>nx38344, A0=>nx38024, A1=>nx38354);
   ix27242 : mux21_ni port map ( Y=>nx27241, A0=>label_4_output_5, A1=>
      label_4_input_5, S0=>nx43431);
   ix12833 : mux21_ni port map ( Y=>nx12832, A0=>nx12828, A1=>
      label_4_input_state_machine_5, S0=>nx42291);
   ix27232 : mux21_ni port map ( Y=>nx27231, A0=>
      label_4_input_state_machine_5, A1=>data_in(53), S0=>nx43381);
   ix38356 : xor2 port map ( Y=>nx38355, A0=>nx38044, A1=>label_4_output_6);
   ix38360 : xnor2 port map ( Y=>nx38359, A0=>nx38063, A1=>nx38369);
   ix27282 : mux21_ni port map ( Y=>nx27281, A0=>label_4_output_7, A1=>
      label_4_input_7, S0=>nx43431);
   ix12897 : mux21_ni port map ( Y=>nx12896, A0=>nx12892, A1=>
      label_4_input_state_machine_7, S0=>nx43085);
   ix27272 : mux21_ni port map ( Y=>nx27271, A0=>
      label_4_input_state_machine_7, A1=>data_in(55), S0=>nx43381);
   ix38371 : xor2 port map ( Y=>nx38370, A0=>nx38096, A1=>label_4_output_8);
   ix38375 : xnor2 port map ( Y=>nx38374, A0=>nx38101, A1=>nx38384);
   ix27322 : mux21_ni port map ( Y=>nx27321, A0=>label_4_output_9, A1=>
      label_4_input_9, S0=>nx43431);
   ix12961 : mux21_ni port map ( Y=>nx12960, A0=>nx12956, A1=>
      label_4_input_state_machine_9, S0=>nx43087);
   ix27312 : mux21_ni port map ( Y=>nx27311, A0=>
      label_4_input_state_machine_9, A1=>data_in(57), S0=>nx43381);
   ix38386 : xor2 port map ( Y=>nx38385, A0=>nx38132, A1=>label_4_output_10
   );
   ix38390 : xnor2 port map ( Y=>nx38389, A0=>nx38137, A1=>nx38399);
   ix27362 : mux21_ni port map ( Y=>nx27361, A0=>label_4_output_11, A1=>
      label_4_input_11, S0=>nx43431);
   ix13025 : mux21_ni port map ( Y=>nx13024, A0=>nx13020, A1=>
      label_4_input_state_machine_11, S0=>nx43087);
   ix27352 : mux21_ni port map ( Y=>nx27351, A0=>
      label_4_input_state_machine_11, A1=>data_in(59), S0=>nx43381);
   ix38401 : xor2 port map ( Y=>nx38400, A0=>nx38168, A1=>label_4_output_12
   );
   ix38405 : xnor2 port map ( Y=>nx38404, A0=>nx38173, A1=>nx38414);
   ix27402 : mux21_ni port map ( Y=>nx27401, A0=>label_4_output_13, A1=>
      label_4_input_13, S0=>nx43431);
   ix13089 : mux21_ni port map ( Y=>nx13088, A0=>nx13084, A1=>
      label_4_input_state_machine_13, S0=>nx43087);
   ix27392 : mux21_ni port map ( Y=>nx27391, A0=>
      label_4_input_state_machine_13, A1=>data_in(61), S0=>nx43381);
   ix38416 : xor2 port map ( Y=>nx38415, A0=>nx38204, A1=>label_4_output_14
   );
   ix16285 : mux21 port map ( Y=>nx16284, A0=>nx39057, A1=>nx38423, S0=>
      nx43013);
   ix28242 : mux21_ni port map ( Y=>nx28241, A0=>label_7_output_14, A1=>
      label_7_input_14, S0=>nx43431);
   ix14425 : mux21_ni port map ( Y=>nx14424, A0=>nx14420, A1=>
      label_7_input_state_machine_14, S0=>nx43087);
   ix27422 : mux21_ni port map ( Y=>nx27421, A0=>
      label_7_input_state_machine_14, A1=>data_in(110), S0=>nx43381);
   ix28212 : mux21_ni port map ( Y=>nx28211, A0=>label_7_output_12, A1=>
      label_7_input_12, S0=>nx43433);
   ix14367 : mux21_ni port map ( Y=>nx14366, A0=>nx14362, A1=>
      label_7_input_state_machine_12, S0=>nx43087);
   ix28202 : mux21_ni port map ( Y=>nx28201, A0=>
      label_7_input_state_machine_12, A1=>data_in(108), S0=>nx43383);
   ix28172 : mux21_ni port map ( Y=>nx28171, A0=>label_7_output_10, A1=>
      label_7_input_10, S0=>nx43433);
   ix14303 : mux21_ni port map ( Y=>nx14302, A0=>nx14298, A1=>
      label_7_input_state_machine_10, S0=>nx43087);
   ix28162 : mux21_ni port map ( Y=>nx28161, A0=>
      label_7_input_state_machine_10, A1=>data_in(106), S0=>nx43383);
   ix28132 : mux21_ni port map ( Y=>nx28131, A0=>label_7_output_8, A1=>
      label_7_input_8, S0=>nx43433);
   ix14239 : mux21_ni port map ( Y=>nx14238, A0=>nx14234, A1=>
      label_7_input_state_machine_8, S0=>nx43087);
   ix28122 : mux21_ni port map ( Y=>nx28121, A0=>
      label_7_input_state_machine_8, A1=>data_in(104), S0=>nx43383);
   ix28092 : mux21_ni port map ( Y=>nx28091, A0=>label_7_output_6, A1=>
      label_7_input_6, S0=>nx43433);
   ix14175 : mux21_ni port map ( Y=>nx14174, A0=>nx14170, A1=>
      label_7_input_state_machine_6, S0=>nx43089);
   ix28082 : mux21_ni port map ( Y=>nx28081, A0=>
      label_7_input_state_machine_6, A1=>data_in(102), S0=>nx43383);
   ix28052 : mux21_ni port map ( Y=>nx28051, A0=>label_7_output_4, A1=>
      label_7_input_4, S0=>nx43433);
   ix14111 : mux21_ni port map ( Y=>nx14110, A0=>nx14106, A1=>
      label_7_input_state_machine_4, S0=>nx43089);
   ix28042 : mux21_ni port map ( Y=>nx28041, A0=>
      label_7_input_state_machine_4, A1=>data_in(100), S0=>nx43383);
   ix28012 : mux21_ni port map ( Y=>nx28011, A0=>label_7_output_2, A1=>
      label_7_input_2, S0=>nx43433);
   ix14047 : mux21_ni port map ( Y=>nx14046, A0=>nx14042, A1=>
      label_7_input_state_machine_2, S0=>nx43089);
   ix28002 : mux21_ni port map ( Y=>nx28001, A0=>
      label_7_input_state_machine_2, A1=>data_in(98), S0=>nx43383);
   ix27972 : mux21_ni port map ( Y=>nx27971, A0=>label_7_output_0, A1=>
      label_7_input_0, S0=>nx43433);
   ix27962 : mux21_ni port map ( Y=>nx27961, A0=>
      label_7_input_state_machine_0, A1=>data_in(96), S0=>nx43383);
   ix27952 : mux21_ni port map ( Y=>nx27951, A0=>
      booth_booth_integration_output_6_12, A1=>nx13966, S0=>nx43305);
   ix13967 : mux21_ni port map ( Y=>nx13966, A0=>nx41809, A1=>
      booth_booth_integration_output_6_13, S0=>nx43313);
   ix27942 : mux21_ni port map ( Y=>nx27941, A0=>
      booth_booth_integration_output_6_13, A1=>nx13954, S0=>nx43305);
   ix13955 : mux21_ni port map ( Y=>nx13954, A0=>nx41805, A1=>
      booth_booth_integration_output_6_14, S0=>nx43313);
   ix27932 : mux21_ni port map ( Y=>nx27931, A0=>
      booth_booth_integration_output_6_14, A1=>nx13942, S0=>nx43305);
   ix13943 : mux21_ni port map ( Y=>nx13942, A0=>nx41801, A1=>
      booth_booth_integration_output_6_15, S0=>nx43313);
   ix27922 : mux21 port map ( Y=>nx27921, A0=>nx38944, A1=>nx38525, S0=>
      nx43305);
   ix27452 : mux21_ni port map ( Y=>nx27451, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_0, A1=>nx42087, S0=>nx42957
   );
   ix27438 : and02 port map ( Y=>nx27437, A0=>nx43495, A1=>
      booth_booth_integrtaion_6_shift_Reg_count_0);
   ix27632 : mux21_ni port map ( Y=>nx27631, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_9, A1=>nx42073, S0=>nx42957
   );
   ix27622 : mux21_ni port map ( Y=>nx27621, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_9, A1=>output_8_dup_12856, 
      S0=>nx43305);
   ix27612 : mux21_ni port map ( Y=>nx27611, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_8, A1=>output_8_dup_12856, 
      S0=>nx42957);
   ix27602 : mux21_ni port map ( Y=>nx27601, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_8, A1=>output_7_dup_12857, 
      S0=>nx43305);
   ix27592 : mux21_ni port map ( Y=>nx27591, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_7, A1=>output_7_dup_12857, 
      S0=>nx42957);
   ix27582 : mux21_ni port map ( Y=>nx27581, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_7, A1=>output_6_dup_12858, 
      S0=>nx43307);
   ix27572 : mux21_ni port map ( Y=>nx27571, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_6, A1=>output_6_dup_12858, 
      S0=>nx42957);
   ix27562 : mux21_ni port map ( Y=>nx27561, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_6, A1=>output_5_dup_12859, 
      S0=>nx43307);
   ix27552 : mux21_ni port map ( Y=>nx27551, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_5, A1=>output_5_dup_12859, 
      S0=>nx42957);
   ix27542 : mux21_ni port map ( Y=>nx27541, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_5, A1=>output_4_dup_12860, 
      S0=>nx43307);
   ix27532 : mux21_ni port map ( Y=>nx27531, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_4, A1=>output_4_dup_12860, 
      S0=>nx42959);
   ix27522 : mux21_ni port map ( Y=>nx27521, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_4, A1=>output_3_dup_12861, 
      S0=>nx43307);
   ix27512 : mux21_ni port map ( Y=>nx27511, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_3, A1=>output_3_dup_12861, 
      S0=>nx42959);
   ix27502 : mux21_ni port map ( Y=>nx27501, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_3, A1=>output_2_dup_12862, 
      S0=>nx43307);
   ix27492 : mux21_ni port map ( Y=>nx27491, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_2, A1=>output_2_dup_12862, 
      S0=>nx42959);
   ix27482 : mux21_ni port map ( Y=>nx27481, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_2, A1=>output_1_dup_12863, 
      S0=>nx43307);
   ix27472 : mux21_ni port map ( Y=>nx27471, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_1, A1=>output_1_dup_12863, 
      S0=>nx42959);
   ix27462 : mux21_ni port map ( Y=>nx27461, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_1, A1=>nx42087, S0=>nx43307
   );
   ix13383 : nand02 port map ( Y=>nx38671, A0=>nx38598, A1=>
      booth_output_0_dup_12225);
   ix38601 : or03 port map ( Y=>nx38600, A0=>nx38649, A1=>
      booth_booth_integrtaion_6_shift_reg_output_0, A2=>nx43495);
   ix27752 : mux21_ni port map ( Y=>nx27751, A0=>booth_output_0_dup_12225, 
      A1=>nx13362, S0=>nx43309);
   ix13363 : mux21_ni port map ( Y=>nx13362, A0=>nx41783, A1=>
      booth_output_1_dup_12224, S0=>nx43315);
   ix27742 : mux21_ni port map ( Y=>nx27741, A0=>booth_output_1_dup_12224, 
      A1=>nx13350, S0=>nx43309);
   ix13351 : mux21_ni port map ( Y=>nx13350, A0=>nx41779, A1=>
      booth_output_2_dup_12223, S0=>nx43315);
   ix27732 : mux21_ni port map ( Y=>nx27731, A0=>booth_output_2_dup_12223, 
      A1=>nx13338, S0=>nx43309);
   ix13339 : mux21_ni port map ( Y=>nx13338, A0=>nx41775, A1=>
      booth_output_3_dup_12222, S0=>nx43315);
   ix27722 : mux21_ni port map ( Y=>nx27721, A0=>booth_output_3_dup_12222, 
      A1=>nx13326, S0=>nx43309);
   ix13327 : mux21_ni port map ( Y=>nx13326, A0=>nx41771, A1=>
      booth_output_4_dup_12221, S0=>nx43315);
   ix27712 : mux21_ni port map ( Y=>nx27711, A0=>booth_output_4_dup_12221, 
      A1=>nx13314, S0=>nx43309);
   ix13315 : mux21_ni port map ( Y=>nx13314, A0=>nx41767, A1=>
      booth_output_5_dup_12220, S0=>nx43315);
   ix27702 : mux21_ni port map ( Y=>nx27701, A0=>booth_output_5_dup_12220, 
      A1=>nx13302, S0=>nx43309);
   ix13303 : mux21_ni port map ( Y=>nx13302, A0=>nx41763, A1=>
      booth_output_6_dup_12219, S0=>nx43315);
   ix27692 : mux21_ni port map ( Y=>nx27691, A0=>booth_output_6_dup_12219, 
      A1=>nx13290, S0=>nx43309);
   ix13291 : mux21_ni port map ( Y=>nx13290, A0=>nx41759, A1=>
      booth_output_7_dup_12218, S0=>nx43315);
   ix27682 : mux21_ni port map ( Y=>nx27681, A0=>booth_output_7_dup_12218, 
      A1=>nx13278, S0=>nx43311);
   ix13279 : mux21_ni port map ( Y=>nx13278, A0=>nx41755, A1=>
      booth_output_8_dup_12217, S0=>nx43317);
   ix27672 : mux21_ni port map ( Y=>nx27671, A0=>booth_output_8_dup_12217, 
      A1=>nx13266, S0=>nx43311);
   ix13267 : mux21_ni port map ( Y=>nx13266, A0=>nx41751, A1=>
      booth_output_9_dup_12216, S0=>nx43317);
   ix27662 : mux21_ni port map ( Y=>nx27661, A0=>booth_output_9_dup_12216, 
      A1=>nx13254, S0=>nx43311);
   ix13255 : mux21_ni port map ( Y=>nx13254, A0=>nx41747, A1=>
      booth_output_10_dup_12215, S0=>nx43317);
   ix27652 : mux21_ni port map ( Y=>nx27651, A0=>booth_output_10_dup_12215, 
      A1=>nx13242, S0=>nx43311);
   ix13243 : mux21_ni port map ( Y=>nx13242, A0=>nx41743, A1=>
      booth_output_11_dup_12214, S0=>nx43317);
   ix27642 : mux21_ni port map ( Y=>nx27641, A0=>booth_output_11_dup_12214, 
      A1=>nx13230, S0=>nx43311);
   ix13231 : mux21_ni port map ( Y=>nx13230, A0=>nx41731, A1=>
      booth_booth_integration_output_6_12, S0=>nx43317);
   ix27912 : mux21_ni port map ( Y=>nx27911, A0=>
      booth_booth_integration_output_6_16, A1=>nx13912, S0=>nx43311);
   ix13913 : nor02ii port map ( Y=>nx13912, A0=>nx38655, A1=>nx43317);
   ix13389 : nor02ii port map ( Y=>nx13388, A0=>nx38593, A1=>
      booth_booth_integration_output_6_16);
   ix13907 : xor2 port map ( Y=>nx18502, A0=>nx38661, A1=>nx38937);
   ix38677 : or02 port map ( Y=>nx38676, A0=>nx38598, A1=>
      booth_output_0_dup_12225);
   ix13895 : xor2 port map ( Y=>nx18503, A0=>nx38681, A1=>nx42735);
   ix38697 : xor2 port map ( Y=>nx38696, A0=>nx38700, A1=>nx13460);
   ix38709 : nor02ii port map ( Y=>nx38708, A0=>nx13426, A1=>data_in(99));
   ix13871 : xor2 port map ( Y=>nx18505, A0=>nx38733, A1=>nx42737);
   ix27872 : mux21_ni port map ( Y=>nx27871, A0=>
      booth_booth_integration_output_6_20, A1=>nx13864, S0=>nx43311);
   ix13865 : nor02ii port map ( Y=>nx13864, A0=>nx38719, A1=>nx43317);
   ix13859 : xor2 port map ( Y=>nx18507, A0=>nx38738, A1=>nx38934);
   ix13847 : xor2 port map ( Y=>nx18508, A0=>nx38769, A1=>nx42739);
   ix27852 : mux21_ni port map ( Y=>nx27851, A0=>
      booth_booth_integration_output_6_22, A1=>nx13840, S0=>nx42729);
   ix13841 : nor02ii port map ( Y=>nx13840, A0=>nx38755, A1=>nx42733);
   ix13835 : xor2 port map ( Y=>nx18509, A0=>nx38774, A1=>nx38931);
   ix13823 : xor2 port map ( Y=>nx18510, A0=>nx38805, A1=>nx42741);
   ix27832 : mux21_ni port map ( Y=>nx27831, A0=>
      booth_booth_integration_output_6_24, A1=>nx13816, S0=>nx42729);
   ix13817 : nor02ii port map ( Y=>nx13816, A0=>nx38791, A1=>nx42733);
   ix13811 : xor2 port map ( Y=>nx18511, A0=>nx38810, A1=>nx38928);
   ix13799 : xor2 port map ( Y=>nx18512, A0=>nx38841, A1=>nx42743);
   ix27812 : mux21_ni port map ( Y=>nx27811, A0=>
      booth_booth_integration_output_6_26, A1=>nx13792, S0=>nx42729);
   ix13793 : nor02ii port map ( Y=>nx13792, A0=>nx38827, A1=>nx42733);
   ix13787 : xor2 port map ( Y=>nx18513, A0=>nx38846, A1=>nx38925);
   ix13775 : xor2 port map ( Y=>nx18515, A0=>nx38877, A1=>nx42745);
   ix27792 : mux21_ni port map ( Y=>nx27791, A0=>booth_output_28_dup_12213, 
      A1=>nx13768, S0=>nx42729);
   ix13769 : nor02ii port map ( Y=>nx13768, A0=>nx38863, A1=>nx42733);
   ix13763 : xor2 port map ( Y=>nx18517, A0=>nx38882, A1=>nx38922);
   ix13751 : xor2 port map ( Y=>nx18519, A0=>nx38898, A1=>nx42747);
   ix38916 : xor2 port map ( Y=>nx38915, A0=>nx38898, A1=>nx13736);
   ix13925 : nor02ii port map ( Y=>nx13924, A0=>nx13388, A1=>nx42733);
   ix38952 : xnor2 port map ( Y=>nx38951, A0=>nx38947, A1=>nx38961);
   ix27992 : mux21_ni port map ( Y=>nx27991, A0=>label_7_output_1, A1=>
      label_7_input_1, S0=>nx43435);
   ix14015 : mux21_ni port map ( Y=>nx14014, A0=>nx14010, A1=>
      label_7_input_state_machine_1, S0=>nx43089);
   ix27982 : mux21_ni port map ( Y=>nx27981, A0=>
      label_7_input_state_machine_1, A1=>data_in(97), S0=>nx42799);
   ix38967 : xnor2 port map ( Y=>nx38966, A0=>nx38944, A1=>nx38976);
   ix28032 : mux21_ni port map ( Y=>nx28031, A0=>label_7_output_3, A1=>
      label_7_input_3, S0=>nx43435);
   ix14079 : mux21_ni port map ( Y=>nx14078, A0=>nx14074, A1=>
      label_7_input_state_machine_3, S0=>nx43089);
   ix28022 : mux21_ni port map ( Y=>nx28021, A0=>
      label_7_input_state_machine_3, A1=>data_in(99), S0=>nx42799);
   ix38978 : xor2 port map ( Y=>nx38977, A0=>nx38651, A1=>label_7_output_4);
   ix38982 : xnor2 port map ( Y=>nx38981, A0=>nx38661, A1=>nx38991);
   ix28072 : mux21_ni port map ( Y=>nx28071, A0=>label_7_output_5, A1=>
      label_7_input_5, S0=>nx43435);
   ix14143 : mux21_ni port map ( Y=>nx14142, A0=>nx14138, A1=>
      label_7_input_state_machine_5, S0=>nx43089);
   ix28062 : mux21_ni port map ( Y=>nx28061, A0=>
      label_7_input_state_machine_5, A1=>data_in(101), S0=>nx42799);
   ix38993 : xor2 port map ( Y=>nx38992, A0=>nx38681, A1=>label_7_output_6);
   ix38997 : xnor2 port map ( Y=>nx38996, A0=>nx38700, A1=>nx39006);
   ix28112 : mux21_ni port map ( Y=>nx28111, A0=>label_7_output_7, A1=>
      label_7_input_7, S0=>nx43435);
   ix14207 : mux21_ni port map ( Y=>nx14206, A0=>nx14202, A1=>
      label_7_input_state_machine_7, S0=>nx43089);
   ix28102 : mux21_ni port map ( Y=>nx28101, A0=>
      label_7_input_state_machine_7, A1=>data_in(103), S0=>nx42799);
   ix39008 : xor2 port map ( Y=>nx39007, A0=>nx38733, A1=>label_7_output_8);
   ix39012 : xnor2 port map ( Y=>nx39011, A0=>nx38738, A1=>nx39021);
   ix28152 : mux21_ni port map ( Y=>nx28151, A0=>label_7_output_9, A1=>
      label_7_input_9, S0=>nx43435);
   ix14271 : mux21_ni port map ( Y=>nx14270, A0=>nx14266, A1=>
      label_7_input_state_machine_9, S0=>nx43091);
   ix28142 : mux21_ni port map ( Y=>nx28141, A0=>
      label_7_input_state_machine_9, A1=>data_in(105), S0=>nx42799);
   ix39023 : xor2 port map ( Y=>nx39022, A0=>nx38769, A1=>label_7_output_10
   );
   ix39027 : xnor2 port map ( Y=>nx39026, A0=>nx38774, A1=>nx39036);
   ix28192 : mux21_ni port map ( Y=>nx28191, A0=>label_7_output_11, A1=>
      label_7_input_11, S0=>nx43435);
   ix14335 : mux21_ni port map ( Y=>nx14334, A0=>nx14330, A1=>
      label_7_input_state_machine_11, S0=>nx43091);
   ix28182 : mux21_ni port map ( Y=>nx28181, A0=>
      label_7_input_state_machine_11, A1=>data_in(107), S0=>nx42799);
   ix39038 : xor2 port map ( Y=>nx39037, A0=>nx38805, A1=>label_7_output_12
   );
   ix39042 : xnor2 port map ( Y=>nx39041, A0=>nx38810, A1=>nx39051);
   ix28232 : mux21_ni port map ( Y=>nx28231, A0=>label_7_output_13, A1=>
      label_7_input_13, S0=>nx43435);
   ix14399 : mux21_ni port map ( Y=>nx14398, A0=>nx14394, A1=>
      label_7_input_state_machine_13, S0=>nx43091);
   ix28222 : mux21_ni port map ( Y=>nx28221, A0=>
      label_7_input_state_machine_13, A1=>data_in(109), S0=>nx42799);
   ix39053 : xor2 port map ( Y=>nx39052, A0=>nx38841, A1=>label_7_output_14
   );
   ix29082 : mux21_ni port map ( Y=>nx29081, A0=>label_8_output_14, A1=>
      label_8_input_14, S0=>nx43437);
   ix15741 : mux21_ni port map ( Y=>nx15740, A0=>nx15736, A1=>
      label_8_input_state_machine_14, S0=>nx43091);
   ix28262 : mux21_ni port map ( Y=>nx28261, A0=>
      label_8_input_state_machine_14, A1=>data_in(126), S0=>nx43385);
   ix29052 : mux21_ni port map ( Y=>nx29051, A0=>label_8_output_12, A1=>
      label_8_input_12, S0=>nx43437);
   ix15683 : mux21_ni port map ( Y=>nx15682, A0=>nx15678, A1=>
      label_8_input_state_machine_12, S0=>nx43091);
   ix29042 : mux21_ni port map ( Y=>nx29041, A0=>
      label_8_input_state_machine_12, A1=>data_in(124), S0=>nx43385);
   ix29012 : mux21_ni port map ( Y=>nx29011, A0=>label_8_output_10, A1=>
      label_8_input_10, S0=>nx43439);
   ix15619 : mux21_ni port map ( Y=>nx15618, A0=>nx15614, A1=>
      label_8_input_state_machine_10, S0=>nx43091);
   ix29002 : mux21_ni port map ( Y=>nx29001, A0=>
      label_8_input_state_machine_10, A1=>data_in(122), S0=>nx43385);
   ix28972 : mux21_ni port map ( Y=>nx28971, A0=>label_8_output_8, A1=>
      label_8_input_8, S0=>nx43439);
   ix15555 : mux21_ni port map ( Y=>nx15554, A0=>nx15550, A1=>
      label_8_input_state_machine_8, S0=>nx43091);
   ix28962 : mux21_ni port map ( Y=>nx28961, A0=>
      label_8_input_state_machine_8, A1=>data_in(120), S0=>nx43385);
   ix28932 : mux21_ni port map ( Y=>nx28931, A0=>label_8_output_6, A1=>
      label_8_input_6, S0=>nx42813);
   ix15491 : mux21_ni port map ( Y=>nx15490, A0=>nx15486, A1=>
      label_8_input_state_machine_6, S0=>nx43093);
   ix28922 : mux21_ni port map ( Y=>nx28921, A0=>
      label_8_input_state_machine_6, A1=>data_in(118), S0=>nx43385);
   ix28892 : mux21_ni port map ( Y=>nx28891, A0=>label_8_output_4, A1=>
      label_8_input_4, S0=>nx42813);
   ix15427 : mux21_ni port map ( Y=>nx15426, A0=>nx15422, A1=>
      label_8_input_state_machine_4, S0=>nx43093);
   ix28882 : mux21_ni port map ( Y=>nx28881, A0=>
      label_8_input_state_machine_4, A1=>data_in(116), S0=>nx43385);
   ix28852 : mux21_ni port map ( Y=>nx28851, A0=>label_8_output_2, A1=>
      label_8_input_2, S0=>nx42813);
   ix15363 : mux21_ni port map ( Y=>nx15362, A0=>nx15358, A1=>
      label_8_input_state_machine_2, S0=>nx43093);
   ix28842 : mux21_ni port map ( Y=>nx28841, A0=>
      label_8_input_state_machine_2, A1=>data_in(114), S0=>nx43385);
   ix28812 : mux21_ni port map ( Y=>nx28811, A0=>label_8_output_0, A1=>
      label_8_input_0, S0=>nx42813);
   ix28802 : mux21_ni port map ( Y=>nx28801, A0=>
      label_8_input_state_machine_0, A1=>data_in(112), S0=>nx43387);
   ix28792 : mux21_ni port map ( Y=>nx28791, A0=>
      booth_booth_integration_output_7_12, A1=>nx15282, S0=>nx43319);
   ix15283 : mux21_ni port map ( Y=>nx15282, A0=>nx41809, A1=>
      booth_booth_integration_output_7_13, S0=>nx43327);
   ix28782 : mux21_ni port map ( Y=>nx28781, A0=>
      booth_booth_integration_output_7_13, A1=>nx15270, S0=>nx43319);
   ix15271 : mux21_ni port map ( Y=>nx15270, A0=>nx41805, A1=>
      booth_booth_integration_output_7_14, S0=>nx43327);
   ix28772 : mux21_ni port map ( Y=>nx28771, A0=>
      booth_booth_integration_output_7_14, A1=>nx15258, S0=>nx43319);
   ix15259 : mux21_ni port map ( Y=>nx15258, A0=>nx41801, A1=>
      booth_booth_integration_output_7_15, S0=>nx43327);
   ix28762 : mux21 port map ( Y=>nx28761, A0=>nx39578, A1=>nx39159, S0=>
      nx43319);
   ix28292 : mux21_ni port map ( Y=>nx28291, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_0, A1=>nx42119, S0=>nx42961
   );
   ix28278 : and02 port map ( Y=>nx28277, A0=>nx43499, A1=>
      booth_booth_integrtaion_7_shift_Reg_count_0);
   ix28472 : mux21_ni port map ( Y=>nx28471, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_9, A1=>nx42105, S0=>nx42961
   );
   ix28462 : mux21_ni port map ( Y=>nx28461, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_9, A1=>output_8_dup_12884, 
      S0=>nx43319);
   ix28452 : mux21_ni port map ( Y=>nx28451, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_8, A1=>output_8_dup_12884, 
      S0=>nx42961);
   ix28442 : mux21_ni port map ( Y=>nx28441, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_8, A1=>output_7_dup_12885, 
      S0=>nx43319);
   ix28432 : mux21_ni port map ( Y=>nx28431, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_7, A1=>output_7_dup_12885, 
      S0=>nx42961);
   ix28422 : mux21_ni port map ( Y=>nx28421, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_7, A1=>output_6_dup_12886, 
      S0=>nx43321);
   ix28412 : mux21_ni port map ( Y=>nx28411, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_6, A1=>output_6_dup_12886, 
      S0=>nx42961);
   ix28402 : mux21_ni port map ( Y=>nx28401, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_6, A1=>output_5_dup_12887, 
      S0=>nx43321);
   ix28392 : mux21_ni port map ( Y=>nx28391, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_5, A1=>output_5_dup_12887, 
      S0=>nx42961);
   ix28382 : mux21_ni port map ( Y=>nx28381, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_5, A1=>output_4_dup_12888, 
      S0=>nx43321);
   ix28372 : mux21_ni port map ( Y=>nx28371, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_4, A1=>output_4_dup_12888, 
      S0=>nx42963);
   ix28362 : mux21_ni port map ( Y=>nx28361, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_4, A1=>output_3_dup_12889, 
      S0=>nx43321);
   ix28352 : mux21_ni port map ( Y=>nx28351, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_3, A1=>output_3_dup_12889, 
      S0=>nx42963);
   ix28342 : mux21_ni port map ( Y=>nx28341, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_3, A1=>output_2_dup_12890, 
      S0=>nx43321);
   ix28332 : mux21_ni port map ( Y=>nx28331, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_2, A1=>output_2_dup_12890, 
      S0=>nx42963);
   ix28322 : mux21_ni port map ( Y=>nx28321, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_2, A1=>output_1_dup_12891, 
      S0=>nx43321);
   ix28312 : mux21_ni port map ( Y=>nx28311, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_1, A1=>output_1_dup_12891, 
      S0=>nx42963);
   ix28302 : mux21_ni port map ( Y=>nx28301, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_1, A1=>nx42119, S0=>nx43321
   );
   ix14699 : nand02 port map ( Y=>nx39305, A0=>nx39232, A1=>
      booth_output_0_dup_12244);
   ix39235 : or03 port map ( Y=>nx39234, A0=>nx39283, A1=>
      booth_booth_integrtaion_7_shift_reg_output_0, A2=>nx43499);
   ix28592 : mux21_ni port map ( Y=>nx28591, A0=>booth_output_0_dup_12244, 
      A1=>nx14678, S0=>nx43323);
   ix14679 : mux21_ni port map ( Y=>nx14678, A0=>nx41783, A1=>
      booth_output_1_dup_12243, S0=>nx43329);
   ix28582 : mux21_ni port map ( Y=>nx28581, A0=>booth_output_1_dup_12243, 
      A1=>nx14666, S0=>nx43323);
   ix14667 : mux21_ni port map ( Y=>nx14666, A0=>nx41779, A1=>
      booth_output_2_dup_12242, S0=>nx43329);
   ix28572 : mux21_ni port map ( Y=>nx28571, A0=>booth_output_2_dup_12242, 
      A1=>nx14654, S0=>nx43323);
   ix14655 : mux21_ni port map ( Y=>nx14654, A0=>nx41775, A1=>
      booth_output_3_dup_12241, S0=>nx43329);
   ix28562 : mux21_ni port map ( Y=>nx28561, A0=>booth_output_3_dup_12241, 
      A1=>nx14642, S0=>nx43323);
   ix14643 : mux21_ni port map ( Y=>nx14642, A0=>nx41771, A1=>
      booth_output_4_dup_12240, S0=>nx43329);
   ix28552 : mux21_ni port map ( Y=>nx28551, A0=>booth_output_4_dup_12240, 
      A1=>nx14630, S0=>nx43323);
   ix14631 : mux21_ni port map ( Y=>nx14630, A0=>nx41767, A1=>
      booth_output_5_dup_12239, S0=>nx43329);
   ix28542 : mux21_ni port map ( Y=>nx28541, A0=>booth_output_5_dup_12239, 
      A1=>nx14618, S0=>nx43323);
   ix14619 : mux21_ni port map ( Y=>nx14618, A0=>nx41763, A1=>
      booth_output_6_dup_12238, S0=>nx43329);
   ix28532 : mux21_ni port map ( Y=>nx28531, A0=>booth_output_6_dup_12238, 
      A1=>nx14606, S0=>nx43323);
   ix14607 : mux21_ni port map ( Y=>nx14606, A0=>nx41759, A1=>
      booth_output_7_dup_12237, S0=>nx43329);
   ix28522 : mux21_ni port map ( Y=>nx28521, A0=>booth_output_7_dup_12237, 
      A1=>nx14594, S0=>nx43325);
   ix14595 : mux21_ni port map ( Y=>nx14594, A0=>nx41755, A1=>
      booth_output_8_dup_12236, S0=>nx43331);
   ix28512 : mux21_ni port map ( Y=>nx28511, A0=>booth_output_8_dup_12236, 
      A1=>nx14582, S0=>nx43325);
   ix14583 : mux21_ni port map ( Y=>nx14582, A0=>nx41751, A1=>
      booth_output_9_dup_12235, S0=>nx43331);
   ix28502 : mux21_ni port map ( Y=>nx28501, A0=>booth_output_9_dup_12235, 
      A1=>nx14570, S0=>nx43325);
   ix14571 : mux21_ni port map ( Y=>nx14570, A0=>nx41747, A1=>
      booth_output_10_dup_12234, S0=>nx43331);
   ix28492 : mux21_ni port map ( Y=>nx28491, A0=>booth_output_10_dup_12234, 
      A1=>nx14558, S0=>nx43325);
   ix14559 : mux21_ni port map ( Y=>nx14558, A0=>nx41743, A1=>
      booth_output_11_dup_12233, S0=>nx43331);
   ix28482 : mux21_ni port map ( Y=>nx28481, A0=>booth_output_11_dup_12233, 
      A1=>nx14546, S0=>nx43325);
   ix14547 : mux21_ni port map ( Y=>nx14546, A0=>nx41731, A1=>
      booth_booth_integration_output_7_12, S0=>nx43331);
   ix28752 : mux21_ni port map ( Y=>nx28751, A0=>
      booth_booth_integration_output_7_16, A1=>nx15228, S0=>nx43325);
   ix15229 : nor02ii port map ( Y=>nx15228, A0=>nx39289, A1=>nx43331);
   ix14705 : nor02ii port map ( Y=>nx14704, A0=>nx39227, A1=>
      booth_booth_integration_output_7_16);
   ix15223 : xor2 port map ( Y=>nx18544, A0=>nx39295, A1=>nx39571);
   ix39311 : or02 port map ( Y=>nx39310, A0=>nx39232, A1=>
      booth_output_0_dup_12244);
   ix15211 : xor2 port map ( Y=>nx18545, A0=>nx39315, A1=>nx42761);
   ix39331 : xor2 port map ( Y=>nx39330, A0=>nx39334, A1=>nx14776);
   ix39343 : nor02ii port map ( Y=>nx39342, A0=>nx14742, A1=>data_in(115));
   ix15187 : xor2 port map ( Y=>nx18547, A0=>nx39367, A1=>nx42763);
   ix28712 : mux21_ni port map ( Y=>nx28711, A0=>
      booth_booth_integration_output_7_20, A1=>nx15180, S0=>nx43325);
   ix15181 : nor02ii port map ( Y=>nx15180, A0=>nx39353, A1=>nx43331);
   ix15175 : xor2 port map ( Y=>nx18548, A0=>nx39372, A1=>nx39568);
   ix15163 : xor2 port map ( Y=>nx18549, A0=>nx39403, A1=>nx42765);
   ix28692 : mux21_ni port map ( Y=>nx28691, A0=>
      booth_booth_integration_output_7_22, A1=>nx15156, S0=>nx42755);
   ix15157 : nor02ii port map ( Y=>nx15156, A0=>nx39389, A1=>nx42759);
   ix15151 : xor2 port map ( Y=>nx18551, A0=>nx39408, A1=>nx39565);
   ix15139 : xor2 port map ( Y=>nx18553, A0=>nx39439, A1=>nx42767);
   ix28672 : mux21_ni port map ( Y=>nx28671, A0=>
      booth_booth_integration_output_7_24, A1=>nx15132, S0=>nx42755);
   ix15133 : nor02ii port map ( Y=>nx15132, A0=>nx39425, A1=>nx42759);
   ix15127 : xor2 port map ( Y=>nx18555, A0=>nx39444, A1=>nx39562);
   ix15115 : xor2 port map ( Y=>nx18557, A0=>nx39475, A1=>nx42769);
   ix28652 : mux21_ni port map ( Y=>nx28651, A0=>
      booth_booth_integration_output_7_26, A1=>nx15108, S0=>nx42755);
   ix15109 : nor02ii port map ( Y=>nx15108, A0=>nx39461, A1=>nx42759);
   ix15103 : xor2 port map ( Y=>nx18559, A0=>nx39480, A1=>nx39559);
   ix15091 : xor2 port map ( Y=>nx18561, A0=>nx39511, A1=>nx42771);
   ix28632 : mux21_ni port map ( Y=>nx28631, A0=>booth_output_28_dup_12232, 
      A1=>nx15084, S0=>nx42755);
   ix15085 : nor02ii port map ( Y=>nx15084, A0=>nx39497, A1=>nx42759);
   ix15079 : xor2 port map ( Y=>nx18562, A0=>nx39516, A1=>nx39556);
   ix15067 : xor2 port map ( Y=>nx18563, A0=>nx39532, A1=>nx42773);
   ix39550 : xor2 port map ( Y=>nx39549, A0=>nx39532, A1=>nx15052);
   ix15241 : nor02ii port map ( Y=>nx15240, A0=>nx14704, A1=>nx42759);
   ix39586 : xnor2 port map ( Y=>nx39585, A0=>nx39581, A1=>nx39595);
   ix28832 : mux21_ni port map ( Y=>nx28831, A0=>label_8_output_1, A1=>
      label_8_input_1, S0=>nx42813);
   ix15331 : mux21_ni port map ( Y=>nx15330, A0=>nx15326, A1=>
      label_8_input_state_machine_1, S0=>nx43093);
   ix28822 : mux21_ni port map ( Y=>nx28821, A0=>
      label_8_input_state_machine_1, A1=>data_in(113), S0=>nx43387);
   ix39601 : xnor2 port map ( Y=>nx39600, A0=>nx39578, A1=>nx39610);
   ix28872 : mux21_ni port map ( Y=>nx28871, A0=>label_8_output_3, A1=>
      label_8_input_3, S0=>nx42813);
   ix15395 : mux21_ni port map ( Y=>nx15394, A0=>nx15390, A1=>
      label_8_input_state_machine_3, S0=>nx43093);
   ix28862 : mux21_ni port map ( Y=>nx28861, A0=>
      label_8_input_state_machine_3, A1=>data_in(115), S0=>nx43387);
   ix39612 : xor2 port map ( Y=>nx39611, A0=>nx39285, A1=>label_8_output_4);
   ix39616 : xnor2 port map ( Y=>nx39615, A0=>nx39295, A1=>nx39625);
   ix28912 : mux21_ni port map ( Y=>nx28911, A0=>label_8_output_5, A1=>
      label_8_input_5, S0=>nx42813);
   ix15459 : mux21_ni port map ( Y=>nx15458, A0=>nx15454, A1=>
      label_8_input_state_machine_5, S0=>nx43093);
   ix28902 : mux21_ni port map ( Y=>nx28901, A0=>
      label_8_input_state_machine_5, A1=>data_in(117), S0=>nx43387);
   ix39627 : xor2 port map ( Y=>nx39626, A0=>nx39315, A1=>label_8_output_6);
   ix39631 : xnor2 port map ( Y=>nx39630, A0=>nx39334, A1=>nx39640);
   ix28952 : mux21_ni port map ( Y=>nx28951, A0=>label_8_output_7, A1=>
      label_8_input_7, S0=>nx43439);
   ix15523 : mux21_ni port map ( Y=>nx15522, A0=>nx15518, A1=>
      label_8_input_state_machine_7, S0=>nx43093);
   ix28942 : mux21_ni port map ( Y=>nx28941, A0=>
      label_8_input_state_machine_7, A1=>data_in(119), S0=>nx43387);
   ix39642 : xor2 port map ( Y=>nx39641, A0=>nx39367, A1=>label_8_output_8);
   ix39646 : xnor2 port map ( Y=>nx39645, A0=>nx39372, A1=>nx39655);
   ix28992 : mux21_ni port map ( Y=>nx28991, A0=>label_8_output_9, A1=>
      label_8_input_9, S0=>nx43439);
   ix15587 : mux21_ni port map ( Y=>nx15586, A0=>nx15582, A1=>
      label_8_input_state_machine_9, S0=>nx43095);
   ix28982 : mux21_ni port map ( Y=>nx28981, A0=>
      label_8_input_state_machine_9, A1=>data_in(121), S0=>nx43387);
   ix39657 : xor2 port map ( Y=>nx39656, A0=>nx39403, A1=>label_8_output_10
   );
   ix39661 : xnor2 port map ( Y=>nx39660, A0=>nx39408, A1=>nx39670);
   ix29032 : mux21_ni port map ( Y=>nx29031, A0=>label_8_output_11, A1=>
      label_8_input_11, S0=>nx43439);
   ix15651 : mux21_ni port map ( Y=>nx15650, A0=>nx15646, A1=>
      label_8_input_state_machine_11, S0=>nx43095);
   ix29022 : mux21_ni port map ( Y=>nx29021, A0=>
      label_8_input_state_machine_11, A1=>data_in(123), S0=>nx43387);
   ix39672 : xor2 port map ( Y=>nx39671, A0=>nx39439, A1=>label_8_output_12
   );
   ix39676 : xnor2 port map ( Y=>nx39675, A0=>nx39444, A1=>nx39685);
   ix29072 : mux21_ni port map ( Y=>nx29071, A0=>label_8_output_13, A1=>
      label_8_input_13, S0=>nx43439);
   ix15715 : mux21_ni port map ( Y=>nx15714, A0=>nx15710, A1=>
      label_8_input_state_machine_13, S0=>nx43095);
   ix29062 : mux21_ni port map ( Y=>nx29061, A0=>
      label_8_input_state_machine_13, A1=>data_in(125), S0=>nx42801);
   ix39687 : xor2 port map ( Y=>nx39686, A0=>nx39475, A1=>label_8_output_14
   );
   ix15763 : xnor2 port map ( Y=>nx15762, A0=>nx39057, A1=>nx38423);
   ix39695 : xnor2 port map ( Y=>nx39694, A0=>nx39698, A1=>
      max_calc_comparator_fourth_inp1_13);
   ix39701 : or03 port map ( Y=>nx39700, A0=>nx39685, A1=>nx43347, A2=>
      nx43215);
   ix39706 : or03 port map ( Y=>nx39705, A0=>nx39051, A1=>nx43263, A2=>
      nx43215);
   ix15807 : xnor2 port map ( Y=>nx15806, A0=>nx39709, A1=>nx39716);
   ix39723 : xnor2 port map ( Y=>nx39722, A0=>nx39726, A1=>
      max_calc_comparator_fourth_inp1_11);
   ix39729 : or03 port map ( Y=>nx39728, A0=>nx39670, A1=>nx43263, A2=>
      nx43215);
   ix39734 : or03 port map ( Y=>nx39733, A0=>nx39036, A1=>nx43263, A2=>
      nx43215);
   ix15851 : xnor2 port map ( Y=>nx15850, A0=>nx39737, A1=>nx39744);
   ix39751 : xnor2 port map ( Y=>nx39750, A0=>nx39754, A1=>
      max_calc_comparator_fourth_inp1_9);
   ix39757 : or03 port map ( Y=>nx39756, A0=>nx39655, A1=>nx43265, A2=>
      nx42545);
   ix39762 : or03 port map ( Y=>nx39761, A0=>nx39021, A1=>nx43265, A2=>
      nx42545);
   ix15895 : xnor2 port map ( Y=>nx15894, A0=>nx39765, A1=>nx39772);
   ix39779 : xnor2 port map ( Y=>nx39778, A0=>nx39782, A1=>
      max_calc_comparator_fourth_inp1_7);
   ix39785 : or03 port map ( Y=>nx39784, A0=>nx39640, A1=>nx43265, A2=>
      nx42545);
   ix39790 : or03 port map ( Y=>nx39789, A0=>nx39006, A1=>nx43265, A2=>
      nx42545);
   ix15939 : xnor2 port map ( Y=>nx15938, A0=>nx39793, A1=>nx39800);
   ix39807 : xnor2 port map ( Y=>nx39806, A0=>nx39810, A1=>
      max_calc_comparator_fourth_inp1_5);
   ix39813 : or03 port map ( Y=>nx39812, A0=>nx39625, A1=>nx43265, A2=>
      nx43219);
   ix39818 : or03 port map ( Y=>nx39817, A0=>nx38991, A1=>nx43265, A2=>
      nx43219);
   ix15983 : xnor2 port map ( Y=>nx15982, A0=>nx39821, A1=>nx39828);
   ix39835 : xnor2 port map ( Y=>nx39834, A0=>nx39838, A1=>
      max_calc_comparator_fourth_inp1_3);
   ix39841 : or03 port map ( Y=>nx39840, A0=>nx39610, A1=>nx43265, A2=>
      nx43219);
   ix39846 : or03 port map ( Y=>nx39845, A0=>nx38976, A1=>nx43267, A2=>
      nx43219);
   ix16027 : xnor2 port map ( Y=>nx16026, A0=>nx39849, A1=>nx39856);
   ix39867 : or03 port map ( Y=>nx39866, A0=>nx39595, A1=>nx43267, A2=>
      nx43219);
   ix39872 : or03 port map ( Y=>nx39871, A0=>nx38961, A1=>nx43267, A2=>
      nx43219);
   ix16049 : xnor2 port map ( Y=>nx16048, A0=>nx39864, A1=>nx39868);
   ix16275 : xnor2 port map ( Y=>nx16274, A0=>nx39890, A1=>nx39910);
   ix39893 : or03 port map ( Y=>nx39892, A0=>nx39906, A1=>nx43267, A2=>
      nx43219);
   ix29392 : mux21_ni port map ( Y=>nx29391, A0=>label_8_output_15, A1=>
      label_8_input_15, S0=>nx43439);
   ix16211 : mux21_ni port map ( Y=>nx16210, A0=>nx16206, A1=>
      label_8_input_state_machine_15, S0=>nx43095);
   ix29382 : mux21_ni port map ( Y=>nx29381, A0=>
      label_8_input_state_machine_15, A1=>data_in(127), S0=>nx42801);
   ix16205 : xnor2 port map ( Y=>nx16204, A0=>nx39480, A1=>label_8_output_15
   );
   ix39913 : or03 port map ( Y=>nx39912, A0=>nx39926, A1=>nx43267, A2=>
      nx42547);
   ix29422 : mux21_ni port map ( Y=>nx29421, A0=>label_7_output_15, A1=>
      label_7_input_15, S0=>nx42815);
   ix16253 : mux21_ni port map ( Y=>nx16252, A0=>nx16248, A1=>
      label_7_input_state_machine_15, S0=>nx43095);
   ix29412 : mux21_ni port map ( Y=>nx29411, A0=>
      label_7_input_state_machine_15, A1=>data_in(111), S0=>nx42801);
   ix16247 : xnor2 port map ( Y=>nx16246, A0=>nx38846, A1=>label_7_output_15
   );
   ix16311 : xnor2 port map ( Y=>nx16310, A0=>nx37785, A1=>nx35633);
   ix39935 : xnor2 port map ( Y=>nx39934, A0=>nx39938, A1=>
      max_calc_comparator_second_inp1_13);
   ix16337 : mux21_ni port map ( Y=>nx16336, A0=>max_calc_ans4_13, A1=>
      label_4_output_13, S0=>nx43139);
   ix16323 : mux21 port map ( Y=>nx16322, A0=>nx39698, A1=>nx39702, S0=>
      nx43013);
   ix16373 : mux21_ni port map ( Y=>nx16372, A0=>max_calc_ans3_13, A1=>
      label_3_output_13, S0=>nx43139);
   ix16359 : mux21 port map ( Y=>nx16358, A0=>nx37548, A1=>nx37552, S0=>
      nx43007);
   ix16411 : mux21_ni port map ( Y=>nx16410, A0=>max_calc_ans4_12, A1=>
      label_4_output_12, S0=>nx43139);
   ix16397 : mux21 port map ( Y=>nx16396, A0=>nx39709, A1=>nx39716, S0=>
      nx43013);
   ix16447 : mux21_ni port map ( Y=>nx16446, A0=>max_calc_ans3_12, A1=>
      label_3_output_12, S0=>nx43139);
   ix16433 : mux21 port map ( Y=>nx16432, A0=>nx37559, A1=>nx37566, S0=>
      nx43007);
   ix16459 : xnor2 port map ( Y=>nx16458, A0=>nx39959, A1=>nx39971);
   ix39983 : xnor2 port map ( Y=>nx39982, A0=>nx39986, A1=>
      max_calc_comparator_second_inp1_11);
   ix16485 : mux21_ni port map ( Y=>nx16484, A0=>max_calc_ans4_11, A1=>
      label_4_output_11, S0=>nx43139);
   ix16471 : mux21 port map ( Y=>nx16470, A0=>nx39726, A1=>nx39730, S0=>
      nx43013);
   ix16521 : mux21_ni port map ( Y=>nx16520, A0=>max_calc_ans3_11, A1=>
      label_3_output_11, S0=>nx43141);
   ix16507 : mux21 port map ( Y=>nx16506, A0=>nx37576, A1=>nx37580, S0=>
      nx43007);
   ix16559 : mux21_ni port map ( Y=>nx16558, A0=>max_calc_ans4_10, A1=>
      label_4_output_10, S0=>nx43141);
   ix16545 : mux21 port map ( Y=>nx16544, A0=>nx39737, A1=>nx39744, S0=>
      nx43013);
   ix16595 : mux21_ni port map ( Y=>nx16594, A0=>max_calc_ans3_10, A1=>
      label_3_output_10, S0=>nx43141);
   ix16581 : mux21 port map ( Y=>nx16580, A0=>nx37587, A1=>nx37594, S0=>
      nx43007);
   ix16607 : xnor2 port map ( Y=>nx16606, A0=>nx40007, A1=>nx40019);
   ix40031 : xnor2 port map ( Y=>nx40030, A0=>nx40034, A1=>
      max_calc_comparator_second_inp1_9);
   ix16633 : mux21_ni port map ( Y=>nx16632, A0=>max_calc_ans4_9, A1=>
      label_4_output_9, S0=>nx43141);
   ix16619 : mux21 port map ( Y=>nx16618, A0=>nx39754, A1=>nx39758, S0=>
      nx43013);
   ix16669 : mux21_ni port map ( Y=>nx16668, A0=>max_calc_ans3_9, A1=>
      label_3_output_9, S0=>nx43141);
   ix16655 : mux21 port map ( Y=>nx16654, A0=>nx37604, A1=>nx37608, S0=>
      nx43007);
   ix16707 : mux21_ni port map ( Y=>nx16706, A0=>max_calc_ans4_8, A1=>
      label_4_output_8, S0=>nx43141);
   ix16693 : mux21 port map ( Y=>nx16692, A0=>nx39765, A1=>nx39772, S0=>
      nx43013);
   ix16743 : mux21_ni port map ( Y=>nx16742, A0=>max_calc_ans3_8, A1=>
      label_3_output_8, S0=>nx43141);
   ix16729 : mux21 port map ( Y=>nx16728, A0=>nx37615, A1=>nx37622, S0=>
      nx43007);
   ix16755 : xnor2 port map ( Y=>nx16754, A0=>nx40055, A1=>nx40067);
   ix40079 : xnor2 port map ( Y=>nx40078, A0=>nx40082, A1=>
      max_calc_comparator_second_inp1_7);
   ix16781 : mux21_ni port map ( Y=>nx16780, A0=>max_calc_ans4_7, A1=>
      label_4_output_7, S0=>nx42453);
   ix16767 : mux21 port map ( Y=>nx16766, A0=>nx39782, A1=>nx39786, S0=>
      nx43015);
   ix16817 : mux21_ni port map ( Y=>nx16816, A0=>max_calc_ans3_7, A1=>
      label_3_output_7, S0=>nx43143);
   ix16803 : mux21 port map ( Y=>nx16802, A0=>nx37632, A1=>nx37636, S0=>
      nx43009);
   ix16855 : mux21_ni port map ( Y=>nx16854, A0=>max_calc_ans4_6, A1=>
      label_4_output_6, S0=>nx43143);
   ix16841 : mux21 port map ( Y=>nx16840, A0=>nx39793, A1=>nx39800, S0=>
      nx43015);
   ix16891 : mux21_ni port map ( Y=>nx16890, A0=>max_calc_ans3_6, A1=>
      label_3_output_6, S0=>nx43143);
   ix16877 : mux21 port map ( Y=>nx16876, A0=>nx37643, A1=>nx37650, S0=>
      nx43009);
   ix16903 : xnor2 port map ( Y=>nx16902, A0=>nx40103, A1=>nx40115);
   ix40127 : xnor2 port map ( Y=>nx40126, A0=>nx40130, A1=>
      max_calc_comparator_second_inp1_5);
   ix16929 : mux21_ni port map ( Y=>nx16928, A0=>max_calc_ans4_5, A1=>
      label_4_output_5, S0=>nx43143);
   ix16915 : mux21 port map ( Y=>nx16914, A0=>nx39810, A1=>nx39814, S0=>
      nx43015);
   ix16965 : mux21_ni port map ( Y=>nx16964, A0=>max_calc_ans3_5, A1=>
      label_3_output_5, S0=>nx43143);
   ix16951 : mux21 port map ( Y=>nx16950, A0=>nx37660, A1=>nx37664, S0=>
      nx43009);
   ix17003 : mux21_ni port map ( Y=>nx17002, A0=>max_calc_ans4_4, A1=>
      label_4_output_4, S0=>nx43143);
   ix16989 : mux21 port map ( Y=>nx16988, A0=>nx39821, A1=>nx39828, S0=>
      nx43015);
   ix17039 : mux21_ni port map ( Y=>nx17038, A0=>max_calc_ans3_4, A1=>
      label_3_output_4, S0=>nx43145);
   ix17025 : mux21 port map ( Y=>nx17024, A0=>nx37671, A1=>nx37678, S0=>
      nx43009);
   ix17051 : xnor2 port map ( Y=>nx17050, A0=>nx40151, A1=>nx40163);
   ix40175 : xnor2 port map ( Y=>nx40174, A0=>nx40178, A1=>
      max_calc_comparator_second_inp1_3);
   ix17077 : mux21_ni port map ( Y=>nx17076, A0=>max_calc_ans4_3, A1=>
      label_4_output_3, S0=>nx43145);
   ix17063 : mux21 port map ( Y=>nx17062, A0=>nx39838, A1=>nx39842, S0=>
      nx43015);
   ix17113 : mux21_ni port map ( Y=>nx17112, A0=>max_calc_ans3_3, A1=>
      label_3_output_3, S0=>nx43145);
   ix17099 : mux21 port map ( Y=>nx17098, A0=>nx37688, A1=>nx37692, S0=>
      nx43009);
   ix17151 : mux21_ni port map ( Y=>nx17150, A0=>max_calc_ans4_2, A1=>
      label_4_output_2, S0=>nx43145);
   ix17137 : mux21 port map ( Y=>nx17136, A0=>nx39849, A1=>nx39856, S0=>
      nx43015);
   ix17187 : mux21_ni port map ( Y=>nx17186, A0=>max_calc_ans3_2, A1=>
      label_3_output_2, S0=>nx43145);
   ix17173 : mux21 port map ( Y=>nx17172, A0=>nx37699, A1=>nx37706, S0=>
      nx43009);
   ix17199 : xnor2 port map ( Y=>nx17198, A0=>nx40199, A1=>nx40211);
   ix17225 : mux21_ni port map ( Y=>nx17224, A0=>max_calc_ans4_1, A1=>
      label_4_output_1, S0=>nx43145);
   ix17211 : mux21 port map ( Y=>nx17210, A0=>nx39864, A1=>nx39868, S0=>
      nx43015);
   ix17261 : mux21_ni port map ( Y=>nx17260, A0=>max_calc_ans3_1, A1=>
      label_3_output_1, S0=>nx43145);
   ix17247 : mux21 port map ( Y=>nx17246, A0=>nx37714, A1=>nx37718, S0=>
      nx43009);
   ix17299 : mux21_ni port map ( Y=>nx17298, A0=>max_calc_ans4_0, A1=>
      label_4_output_0, S0=>nx43147);
   ix17285 : mux21 port map ( Y=>nx17284, A0=>nx39875, A1=>nx39882, S0=>
      nx43017);
   ix17335 : mux21_ni port map ( Y=>nx17334, A0=>max_calc_ans3_0, A1=>
      label_3_output_0, S0=>nx43147);
   ix17321 : mux21 port map ( Y=>nx17320, A0=>nx37725, A1=>nx37732, S0=>
      nx43011);
   ix17273 : xnor2 port map ( Y=>nx17272, A0=>nx40224, A1=>nx40233);
   ix17603 : xnor2 port map ( Y=>nx17602, A0=>nx40270, A1=>nx40295);
   ix17523 : mux21_ni port map ( Y=>nx17522, A0=>max_calc_ans4_15, A1=>
      label_4_output_15, S0=>nx43147);
   ix30032 : mux21_ni port map ( Y=>nx30031, A0=>label_4_output_15, A1=>
      label_4_input_15, S0=>nx42815);
   ix17487 : mux21_ni port map ( Y=>nx17486, A0=>nx17482, A1=>
      label_4_input_state_machine_15, S0=>nx43095);
   ix30022 : mux21_ni port map ( Y=>nx30021, A0=>
      label_4_input_state_machine_15, A1=>data_in(63), S0=>nx42801);
   ix17481 : xnor2 port map ( Y=>nx17480, A0=>nx38209, A1=>label_4_output_15
   );
   ix17509 : mux21 port map ( Y=>nx17508, A0=>nx39890, A1=>nx39910, S0=>
      nx43017);
   ix17591 : mux21_ni port map ( Y=>nx17590, A0=>max_calc_ans3_15, A1=>
      label_3_output_15, S0=>nx43147);
   ix30072 : mux21_ni port map ( Y=>nx30071, A0=>label_3_output_15, A1=>
      label_3_input_15, S0=>nx42815);
   ix17555 : mux21_ni port map ( Y=>nx17554, A0=>nx17550, A1=>
      label_3_input_state_machine_15, S0=>nx43095);
   ix30062 : mux21_ni port map ( Y=>nx30061, A0=>
      label_3_input_state_machine_15, A1=>data_in(47), S0=>nx42801);
   ix17549 : xnor2 port map ( Y=>nx17548, A0=>nx36057, A1=>label_3_output_15
   );
   ix17577 : mux21 port map ( Y=>nx17576, A0=>nx37740, A1=>nx37760, S0=>
      nx43011);
   ix18153 : mux21_ni port map ( Y=>nx18152, A0=>max_calc_ans8_14, A1=>
      max_calc_ans7_14, S0=>nx43147);
   ix30442 : mux21_ni port map ( Y=>nx30441, A0=>max_calc_ans7_14, A1=>
      nx17612, S0=>nx43179);
   ix30432 : mux21_ni port map ( Y=>nx30431, A0=>max_calc_ans8_14, A1=>
      nx18603, S0=>nx43285);
   ix18165 : xor2 port map ( Y=>nx18164, A0=>nx40326, A1=>
      max_calc_comparator_first_inp1_14);
   ix40333 : xor2 port map ( Y=>nx40332, A0=>
      max_calc_comparator_first_inp2_13, A1=>
      max_calc_comparator_first_inp1_13);
   ix30532 : mux21_ni port map ( Y=>nx30531, A0=>
      max_calc_comparator_first_inp2_13, A1=>nx18278, S0=>nx43391);
   ix18279 : mux21_ni port map ( Y=>nx18278, A0=>nx18274, A1=>nx18186, S0=>
      nx43031);
   ix18187 : mux21_ni port map ( Y=>nx18186, A0=>max_calc_ans2_13, A1=>
      label_2_output_13, S0=>nx43147);
   ix30462 : mux21_ni port map ( Y=>nx30461, A0=>nx18176, A1=>
      max_calc_ans2_13, S0=>nx42991);
   ix18177 : mux21 port map ( Y=>nx18176, A0=>nx39938, A1=>nx39947, S0=>
      nx43019);
   ix18275 : mux21_ni port map ( Y=>nx18274, A0=>max_calc_ans8_13, A1=>
      max_calc_ans7_13, S0=>nx43147);
   ix30522 : mux21_ni port map ( Y=>nx30521, A0=>max_calc_ans7_13, A1=>
      nx18176, S0=>nx43179);
   ix30512 : mux21_ni port map ( Y=>nx30511, A0=>max_calc_ans8_13, A1=>
      nx18607, S0=>nx43285);
   ix18255 : mux21_ni port map ( Y=>nx18607, A0=>
      max_calc_comparator_first_inp2_13, A1=>
      max_calc_comparator_first_inp1_13, S0=>nx43025);
   ix30502 : mux21_ni port map ( Y=>nx30501, A0=>
      max_calc_comparator_first_inp1_13, A1=>nx18240, S0=>nx43391);
   ix18241 : mux21_ni port map ( Y=>nx18240, A0=>nx18236, A1=>nx18204, S0=>
      nx43033);
   ix18205 : mux21_ni port map ( Y=>nx18204, A0=>max_calc_ans1_13, A1=>
      label_1_output_13, S0=>nx43149);
   ix30472 : mux21_ni port map ( Y=>nx30471, A0=>nx18607, A1=>
      max_calc_ans1_13, S0=>nx42991);
   ix18237 : mux21_ni port map ( Y=>nx18236, A0=>max_calc_ans5_13, A1=>
      max_calc_ans6_13, S0=>nx43149);
   ix30482 : mux21_ni port map ( Y=>nx30481, A0=>max_calc_ans6_13, A1=>
      nx18607, S0=>nx43179);
   ix30492 : mux21_ni port map ( Y=>nx30491, A0=>max_calc_ans5_13, A1=>
      nx18226, S0=>nx42871);
   ix18227 : mux21 port map ( Y=>nx18226, A0=>nx34773, A1=>nx34777, S0=>
      nx43001);
   ix30612 : mux21_ni port map ( Y=>nx30611, A0=>
      max_calc_comparator_first_inp2_12, A1=>nx18400, S0=>nx43391);
   ix18401 : mux21_ni port map ( Y=>nx18400, A0=>nx18396, A1=>nx18308, S0=>
      nx43033);
   ix18309 : mux21_ni port map ( Y=>nx18308, A0=>max_calc_ans2_12, A1=>
      label_2_output_12, S0=>nx43149);
   ix30542 : mux21_ni port map ( Y=>nx30541, A0=>nx18298, A1=>
      max_calc_ans2_12, S0=>nx42991);
   ix18299 : mux21 port map ( Y=>nx18298, A0=>nx39959, A1=>nx39971, S0=>
      nx43019);
   ix18397 : mux21_ni port map ( Y=>nx18396, A0=>max_calc_ans8_12, A1=>
      max_calc_ans7_12, S0=>nx43149);
   ix30602 : mux21_ni port map ( Y=>nx30601, A0=>max_calc_ans7_12, A1=>
      nx18298, S0=>nx43179);
   ix30592 : mux21_ni port map ( Y=>nx30591, A0=>max_calc_ans8_12, A1=>
      nx18608, S0=>nx43285);
   ix18377 : mux21_ni port map ( Y=>nx18608, A0=>
      max_calc_comparator_first_inp2_12, A1=>
      max_calc_comparator_first_inp1_12, S0=>nx43025);
   ix30582 : mux21_ni port map ( Y=>nx30581, A0=>
      max_calc_comparator_first_inp1_12, A1=>nx18362, S0=>nx43393);
   ix18363 : mux21_ni port map ( Y=>nx18362, A0=>nx18358, A1=>nx18326, S0=>
      nx43033);
   ix18327 : mux21_ni port map ( Y=>nx18326, A0=>max_calc_ans1_12, A1=>
      label_1_output_12, S0=>nx43149);
   ix30552 : mux21_ni port map ( Y=>nx30551, A0=>nx18608, A1=>
      max_calc_ans1_12, S0=>nx42991);
   ix18359 : mux21_ni port map ( Y=>nx18358, A0=>max_calc_ans5_12, A1=>
      max_calc_ans6_12, S0=>nx43149);
   ix30562 : mux21_ni port map ( Y=>nx30561, A0=>max_calc_ans6_12, A1=>
      nx18608, S0=>nx43179);
   ix30572 : mux21_ni port map ( Y=>nx30571, A0=>max_calc_ans5_12, A1=>
      nx18348, S0=>nx42871);
   ix18349 : mux21 port map ( Y=>nx18348, A0=>nx34784, A1=>nx34791, S0=>
      nx43001);
   ix18409 : xor2 port map ( Y=>nx18408, A0=>nx40369, A1=>
      max_calc_comparator_first_inp1_12);
   ix40406 : xor2 port map ( Y=>nx40405, A0=>
      max_calc_comparator_first_inp2_11, A1=>
      max_calc_comparator_first_inp1_11);
   ix30692 : mux21_ni port map ( Y=>nx30691, A0=>
      max_calc_comparator_first_inp2_11, A1=>nx18522, S0=>nx43393);
   ix18523 : mux21_ni port map ( Y=>nx18522, A0=>nx18518, A1=>nx18430, S0=>
      nx43033);
   ix18431 : mux21_ni port map ( Y=>nx18430, A0=>max_calc_ans2_11, A1=>
      label_2_output_11, S0=>nx43149);
   ix30622 : mux21_ni port map ( Y=>nx30621, A0=>nx18420, A1=>
      max_calc_ans2_11, S0=>nx42993);
   ix18421 : mux21 port map ( Y=>nx18420, A0=>nx39986, A1=>nx39995, S0=>
      nx43019);
   ix18519 : mux21_ni port map ( Y=>nx18518, A0=>max_calc_ans8_11, A1=>
      max_calc_ans7_11, S0=>nx43151);
   ix30682 : mux21_ni port map ( Y=>nx30681, A0=>max_calc_ans7_11, A1=>
      nx18420, S0=>nx43179);
   ix30672 : mux21_ni port map ( Y=>nx30671, A0=>max_calc_ans8_11, A1=>
      nx18609, S0=>nx43285);
   ix18499 : mux21_ni port map ( Y=>nx18609, A0=>
      max_calc_comparator_first_inp2_11, A1=>
      max_calc_comparator_first_inp1_11, S0=>nx43025);
   ix30662 : mux21_ni port map ( Y=>nx30661, A0=>
      max_calc_comparator_first_inp1_11, A1=>nx18484, S0=>nx43393);
   ix18485 : mux21_ni port map ( Y=>nx18484, A0=>nx18480, A1=>nx18448, S0=>
      nx43033);
   ix18449 : mux21_ni port map ( Y=>nx18448, A0=>max_calc_ans1_11, A1=>
      label_1_output_11, S0=>nx43151);
   ix30632 : mux21_ni port map ( Y=>nx30631, A0=>nx18609, A1=>
      max_calc_ans1_11, S0=>nx42993);
   ix18481 : mux21_ni port map ( Y=>nx18480, A0=>max_calc_ans5_11, A1=>
      max_calc_ans6_11, S0=>nx43151);
   ix30642 : mux21_ni port map ( Y=>nx30641, A0=>max_calc_ans6_11, A1=>
      nx18609, S0=>nx43181);
   ix30652 : mux21_ni port map ( Y=>nx30651, A0=>max_calc_ans5_11, A1=>
      nx18470, S0=>nx42871);
   ix18471 : mux21 port map ( Y=>nx18470, A0=>nx34801, A1=>nx34805, S0=>
      nx43001);
   ix30772 : mux21_ni port map ( Y=>nx30771, A0=>
      max_calc_comparator_first_inp2_10, A1=>nx18644, S0=>nx43393);
   ix18645 : mux21_ni port map ( Y=>nx18644, A0=>nx18640, A1=>nx18552, S0=>
      nx43033);
   ix18553 : mux21_ni port map ( Y=>nx18552, A0=>max_calc_ans2_10, A1=>
      label_2_output_10, S0=>nx43151);
   ix30702 : mux21_ni port map ( Y=>nx30701, A0=>nx18542, A1=>
      max_calc_ans2_10, S0=>nx42993);
   ix18543 : mux21 port map ( Y=>nx18542, A0=>nx40007, A1=>nx40019, S0=>
      nx43019);
   ix18641 : mux21_ni port map ( Y=>nx18640, A0=>max_calc_ans8_10, A1=>
      max_calc_ans7_10, S0=>nx43151);
   ix30762 : mux21_ni port map ( Y=>nx30761, A0=>max_calc_ans7_10, A1=>
      nx18542, S0=>nx43181);
   ix30752 : mux21_ni port map ( Y=>nx30751, A0=>max_calc_ans8_10, A1=>
      nx18610, S0=>nx43285);
   ix18621 : mux21_ni port map ( Y=>nx18610, A0=>
      max_calc_comparator_first_inp2_10, A1=>
      max_calc_comparator_first_inp1_10, S0=>nx43025);
   ix30742 : mux21_ni port map ( Y=>nx30741, A0=>
      max_calc_comparator_first_inp1_10, A1=>nx18606, S0=>nx43393);
   ix18607 : mux21_ni port map ( Y=>nx18606, A0=>nx18602, A1=>nx18570, S0=>
      nx43033);
   ix18571 : mux21_ni port map ( Y=>nx18570, A0=>max_calc_ans1_10, A1=>
      label_1_output_10, S0=>nx43151);
   ix30712 : mux21_ni port map ( Y=>nx30711, A0=>nx18610, A1=>
      max_calc_ans1_10, S0=>nx42993);
   ix18603 : mux21_ni port map ( Y=>nx18602, A0=>max_calc_ans5_10, A1=>
      max_calc_ans6_10, S0=>nx43151);
   ix30722 : mux21_ni port map ( Y=>nx30721, A0=>max_calc_ans6_10, A1=>
      nx18610, S0=>nx43181);
   ix30732 : mux21_ni port map ( Y=>nx30731, A0=>max_calc_ans5_10, A1=>
      nx18592, S0=>nx42871);
   ix18593 : mux21 port map ( Y=>nx18592, A0=>nx34812, A1=>nx34819, S0=>
      nx43001);
   ix18653 : xor2 port map ( Y=>nx18652, A0=>nx40442, A1=>
      max_calc_comparator_first_inp1_10);
   ix40479 : xor2 port map ( Y=>nx40478, A0=>
      max_calc_comparator_first_inp2_9, A1=>max_calc_comparator_first_inp1_9
   );
   ix30852 : mux21_ni port map ( Y=>nx30851, A0=>
      max_calc_comparator_first_inp2_9, A1=>nx18766, S0=>nx43393);
   ix18767 : mux21_ni port map ( Y=>nx18766, A0=>nx18762, A1=>nx18674, S0=>
      nx43035);
   ix18675 : mux21_ni port map ( Y=>nx18674, A0=>max_calc_ans2_9, A1=>
      label_2_output_9, S0=>nx43153);
   ix30782 : mux21_ni port map ( Y=>nx30781, A0=>nx18664, A1=>
      max_calc_ans2_9, S0=>nx42993);
   ix18665 : mux21 port map ( Y=>nx18664, A0=>nx40034, A1=>nx40043, S0=>
      nx43019);
   ix18763 : mux21_ni port map ( Y=>nx18762, A0=>max_calc_ans8_9, A1=>
      max_calc_ans7_9, S0=>nx43153);
   ix30842 : mux21_ni port map ( Y=>nx30841, A0=>max_calc_ans7_9, A1=>
      nx18664, S0=>nx43181);
   ix30832 : mux21_ni port map ( Y=>nx30831, A0=>max_calc_ans8_9, A1=>
      nx18611, S0=>nx43285);
   ix18743 : mux21_ni port map ( Y=>nx18611, A0=>
      max_calc_comparator_first_inp2_9, A1=>max_calc_comparator_first_inp1_9, 
      S0=>nx43025);
   ix30822 : mux21_ni port map ( Y=>nx30821, A0=>
      max_calc_comparator_first_inp1_9, A1=>nx18728, S0=>nx43393);
   ix18729 : mux21_ni port map ( Y=>nx18728, A0=>nx18724, A1=>nx18692, S0=>
      nx43035);
   ix18693 : mux21_ni port map ( Y=>nx18692, A0=>max_calc_ans1_9, A1=>
      label_1_output_9, S0=>nx43153);
   ix30792 : mux21_ni port map ( Y=>nx30791, A0=>nx18611, A1=>
      max_calc_ans1_9, S0=>nx42993);
   ix18725 : mux21_ni port map ( Y=>nx18724, A0=>max_calc_ans5_9, A1=>
      max_calc_ans6_9, S0=>nx43153);
   ix30802 : mux21_ni port map ( Y=>nx30801, A0=>max_calc_ans6_9, A1=>
      nx18611, S0=>nx43181);
   ix30812 : mux21_ni port map ( Y=>nx30811, A0=>max_calc_ans5_9, A1=>
      nx18714, S0=>nx42873);
   ix18715 : mux21 port map ( Y=>nx18714, A0=>nx34829, A1=>nx34833, S0=>
      nx43001);
   ix30932 : mux21_ni port map ( Y=>nx30931, A0=>
      max_calc_comparator_first_inp2_8, A1=>nx18888, S0=>nx43395);
   ix18889 : mux21_ni port map ( Y=>nx18888, A0=>nx18884, A1=>nx18796, S0=>
      nx43035);
   ix18797 : mux21_ni port map ( Y=>nx18796, A0=>max_calc_ans2_8, A1=>
      label_2_output_8, S0=>nx43153);
   ix30862 : mux21_ni port map ( Y=>nx30861, A0=>nx18786, A1=>
      max_calc_ans2_8, S0=>nx42993);
   ix18787 : mux21 port map ( Y=>nx18786, A0=>nx40055, A1=>nx40067, S0=>
      nx43019);
   ix18885 : mux21_ni port map ( Y=>nx18884, A0=>max_calc_ans8_8, A1=>
      max_calc_ans7_8, S0=>nx43153);
   ix30922 : mux21_ni port map ( Y=>nx30921, A0=>max_calc_ans7_8, A1=>
      nx18786, S0=>nx43181);
   ix30912 : mux21_ni port map ( Y=>nx30911, A0=>max_calc_ans8_8, A1=>
      nx18612, S0=>nx43287);
   ix18865 : mux21_ni port map ( Y=>nx18612, A0=>
      max_calc_comparator_first_inp2_8, A1=>max_calc_comparator_first_inp1_8, 
      S0=>nx43027);
   ix30902 : mux21_ni port map ( Y=>nx30901, A0=>
      max_calc_comparator_first_inp1_8, A1=>nx18850, S0=>nx43395);
   ix18851 : mux21_ni port map ( Y=>nx18850, A0=>nx18846, A1=>nx18814, S0=>
      nx43035);
   ix18815 : mux21_ni port map ( Y=>nx18814, A0=>max_calc_ans1_8, A1=>
      label_1_output_8, S0=>nx43153);
   ix30872 : mux21_ni port map ( Y=>nx30871, A0=>nx18612, A1=>
      max_calc_ans1_8, S0=>nx42995);
   ix18847 : mux21_ni port map ( Y=>nx18846, A0=>max_calc_ans5_8, A1=>
      max_calc_ans6_8, S0=>nx42455);
   ix30882 : mux21_ni port map ( Y=>nx30881, A0=>max_calc_ans6_8, A1=>
      nx18612, S0=>nx43181);
   ix30892 : mux21_ni port map ( Y=>nx30891, A0=>max_calc_ans5_8, A1=>
      nx18836, S0=>nx42873);
   ix18837 : mux21 port map ( Y=>nx18836, A0=>nx34840, A1=>nx34847, S0=>
      nx43001);
   ix18897 : xor2 port map ( Y=>nx18896, A0=>nx40515, A1=>
      max_calc_comparator_first_inp1_8);
   ix40552 : xor2 port map ( Y=>nx40551, A0=>
      max_calc_comparator_first_inp2_7, A1=>max_calc_comparator_first_inp1_7
   );
   ix31012 : mux21_ni port map ( Y=>nx31011, A0=>
      max_calc_comparator_first_inp2_7, A1=>nx19010, S0=>nx43395);
   ix19011 : mux21_ni port map ( Y=>nx19010, A0=>nx19006, A1=>nx18918, S0=>
      nx43035);
   ix18919 : mux21_ni port map ( Y=>nx18918, A0=>max_calc_ans2_7, A1=>
      label_2_output_7, S0=>nx42455);
   ix30942 : mux21_ni port map ( Y=>nx30941, A0=>nx18908, A1=>
      max_calc_ans2_7, S0=>nx42995);
   ix18909 : mux21 port map ( Y=>nx18908, A0=>nx40082, A1=>nx40091, S0=>
      nx43021);
   ix19007 : mux21_ni port map ( Y=>nx19006, A0=>max_calc_ans8_7, A1=>
      max_calc_ans7_7, S0=>nx42455);
   ix31002 : mux21_ni port map ( Y=>nx31001, A0=>max_calc_ans7_7, A1=>
      nx18908, S0=>nx43183);
   ix30992 : mux21_ni port map ( Y=>nx30991, A0=>max_calc_ans8_7, A1=>
      nx18613, S0=>nx43287);
   ix18987 : mux21_ni port map ( Y=>nx18613, A0=>
      max_calc_comparator_first_inp2_7, A1=>max_calc_comparator_first_inp1_7, 
      S0=>nx43027);
   ix30982 : mux21_ni port map ( Y=>nx30981, A0=>
      max_calc_comparator_first_inp1_7, A1=>nx18972, S0=>nx43395);
   ix18973 : mux21_ni port map ( Y=>nx18972, A0=>nx18968, A1=>nx18936, S0=>
      nx43035);
   ix18937 : mux21_ni port map ( Y=>nx18936, A0=>max_calc_ans1_7, A1=>
      label_1_output_7, S0=>nx42455);
   ix30952 : mux21_ni port map ( Y=>nx30951, A0=>nx18613, A1=>
      max_calc_ans1_7, S0=>nx42995);
   ix18969 : mux21_ni port map ( Y=>nx18968, A0=>max_calc_ans5_7, A1=>
      max_calc_ans6_7, S0=>nx42455);
   ix30962 : mux21_ni port map ( Y=>nx30961, A0=>max_calc_ans6_7, A1=>
      nx18613, S0=>nx43183);
   ix30972 : mux21_ni port map ( Y=>nx30971, A0=>max_calc_ans5_7, A1=>
      nx18958, S0=>nx42873);
   ix18959 : mux21 port map ( Y=>nx18958, A0=>nx34857, A1=>nx34861, S0=>
      nx43003);
   ix31092 : mux21_ni port map ( Y=>nx31091, A0=>
      max_calc_comparator_first_inp2_6, A1=>nx19132, S0=>nx43395);
   ix19133 : mux21_ni port map ( Y=>nx19132, A0=>nx19128, A1=>nx19040, S0=>
      nx43035);
   ix19041 : mux21_ni port map ( Y=>nx19040, A0=>max_calc_ans2_6, A1=>
      label_2_output_6, S0=>nx42455);
   ix31022 : mux21_ni port map ( Y=>nx31021, A0=>nx19030, A1=>
      max_calc_ans2_6, S0=>nx42995);
   ix19031 : mux21 port map ( Y=>nx19030, A0=>nx40103, A1=>nx40115, S0=>
      nx43021);
   ix19129 : mux21_ni port map ( Y=>nx19128, A0=>max_calc_ans8_6, A1=>
      max_calc_ans7_6, S0=>nx43155);
   ix31082 : mux21_ni port map ( Y=>nx31081, A0=>max_calc_ans7_6, A1=>
      nx19030, S0=>nx43183);
   ix31072 : mux21_ni port map ( Y=>nx31071, A0=>max_calc_ans8_6, A1=>
      nx18615, S0=>nx43287);
   ix19109 : mux21_ni port map ( Y=>nx18615, A0=>
      max_calc_comparator_first_inp2_6, A1=>max_calc_comparator_first_inp1_6, 
      S0=>nx43027);
   ix31062 : mux21_ni port map ( Y=>nx31061, A0=>
      max_calc_comparator_first_inp1_6, A1=>nx19094, S0=>nx43395);
   ix19095 : mux21_ni port map ( Y=>nx19094, A0=>nx19090, A1=>nx19058, S0=>
      nx43037);
   ix19059 : mux21_ni port map ( Y=>nx19058, A0=>max_calc_ans1_6, A1=>
      label_1_output_6, S0=>nx42455);
   ix31032 : mux21_ni port map ( Y=>nx31031, A0=>nx18615, A1=>
      max_calc_ans1_6, S0=>nx42995);
   ix19091 : mux21_ni port map ( Y=>nx19090, A0=>max_calc_ans5_6, A1=>
      max_calc_ans6_6, S0=>nx43155);
   ix31042 : mux21_ni port map ( Y=>nx31041, A0=>max_calc_ans6_6, A1=>
      nx18615, S0=>nx43183);
   ix31052 : mux21_ni port map ( Y=>nx31051, A0=>max_calc_ans5_6, A1=>
      nx19080, S0=>nx42873);
   ix19081 : mux21 port map ( Y=>nx19080, A0=>nx34868, A1=>nx34875, S0=>
      nx43003);
   ix19141 : xor2 port map ( Y=>nx19140, A0=>nx40588, A1=>
      max_calc_comparator_first_inp1_6);
   ix40625 : xor2 port map ( Y=>nx40624, A0=>
      max_calc_comparator_first_inp2_5, A1=>max_calc_comparator_first_inp1_5
   );
   ix31172 : mux21_ni port map ( Y=>nx31171, A0=>
      max_calc_comparator_first_inp2_5, A1=>nx19254, S0=>nx43395);
   ix19255 : mux21_ni port map ( Y=>nx19254, A0=>nx19250, A1=>nx19162, S0=>
      nx43037);
   ix19163 : mux21_ni port map ( Y=>nx19162, A0=>max_calc_ans2_5, A1=>
      label_2_output_5, S0=>nx43155);
   ix31102 : mux21_ni port map ( Y=>nx31101, A0=>nx19152, A1=>
      max_calc_ans2_5, S0=>nx42995);
   ix19153 : mux21 port map ( Y=>nx19152, A0=>nx40130, A1=>nx40139, S0=>
      nx43021);
   ix19251 : mux21_ni port map ( Y=>nx19250, A0=>max_calc_ans8_5, A1=>
      max_calc_ans7_5, S0=>nx43155);
   ix31162 : mux21_ni port map ( Y=>nx31161, A0=>max_calc_ans7_5, A1=>
      nx19152, S0=>nx43183);
   ix31152 : mux21_ni port map ( Y=>nx31151, A0=>max_calc_ans8_5, A1=>
      nx18617, S0=>nx43287);
   ix19231 : mux21_ni port map ( Y=>nx18617, A0=>
      max_calc_comparator_first_inp2_5, A1=>max_calc_comparator_first_inp1_5, 
      S0=>nx43027);
   ix31142 : mux21_ni port map ( Y=>nx31141, A0=>
      max_calc_comparator_first_inp1_5, A1=>nx19216, S0=>nx43397);
   ix19217 : mux21_ni port map ( Y=>nx19216, A0=>nx19212, A1=>nx19180, S0=>
      nx43037);
   ix19181 : mux21_ni port map ( Y=>nx19180, A0=>max_calc_ans1_5, A1=>
      label_1_output_5, S0=>nx43155);
   ix31112 : mux21_ni port map ( Y=>nx31111, A0=>nx18617, A1=>
      max_calc_ans1_5, S0=>nx42995);
   ix19213 : mux21_ni port map ( Y=>nx19212, A0=>max_calc_ans5_5, A1=>
      max_calc_ans6_5, S0=>nx43157);
   ix31122 : mux21_ni port map ( Y=>nx31121, A0=>max_calc_ans6_5, A1=>
      nx18617, S0=>nx43183);
   ix31132 : mux21_ni port map ( Y=>nx31131, A0=>max_calc_ans5_5, A1=>
      nx19202, S0=>nx42873);
   ix19203 : mux21 port map ( Y=>nx19202, A0=>nx34885, A1=>nx34889, S0=>
      nx43003);
   ix31252 : mux21_ni port map ( Y=>nx31251, A0=>
      max_calc_comparator_first_inp2_4, A1=>nx19376, S0=>nx43397);
   ix19377 : mux21_ni port map ( Y=>nx19376, A0=>nx19372, A1=>nx19284, S0=>
      nx43037);
   ix19285 : mux21_ni port map ( Y=>nx19284, A0=>max_calc_ans2_4, A1=>
      label_2_output_4, S0=>nx43157);
   ix31182 : mux21_ni port map ( Y=>nx31181, A0=>nx19274, A1=>
      max_calc_ans2_4, S0=>nx42997);
   ix19275 : mux21 port map ( Y=>nx19274, A0=>nx40151, A1=>nx40163, S0=>
      nx43021);
   ix19373 : mux21_ni port map ( Y=>nx19372, A0=>max_calc_ans8_4, A1=>
      max_calc_ans7_4, S0=>nx43157);
   ix31242 : mux21_ni port map ( Y=>nx31241, A0=>max_calc_ans7_4, A1=>
      nx19274, S0=>nx43183);
   ix31232 : mux21_ni port map ( Y=>nx31231, A0=>max_calc_ans8_4, A1=>
      nx18619, S0=>nx43287);
   ix19353 : mux21_ni port map ( Y=>nx18619, A0=>
      max_calc_comparator_first_inp2_4, A1=>max_calc_comparator_first_inp1_4, 
      S0=>nx43027);
   ix31222 : mux21_ni port map ( Y=>nx31221, A0=>
      max_calc_comparator_first_inp1_4, A1=>nx19338, S0=>nx43397);
   ix19339 : mux21_ni port map ( Y=>nx19338, A0=>nx19334, A1=>nx19302, S0=>
      nx43037);
   ix19303 : mux21_ni port map ( Y=>nx19302, A0=>max_calc_ans1_4, A1=>
      label_1_output_4, S0=>nx43157);
   ix31192 : mux21_ni port map ( Y=>nx31191, A0=>nx18619, A1=>
      max_calc_ans1_4, S0=>nx42997);
   ix19335 : mux21_ni port map ( Y=>nx19334, A0=>max_calc_ans5_4, A1=>
      max_calc_ans6_4, S0=>nx43157);
   ix31202 : mux21_ni port map ( Y=>nx31201, A0=>max_calc_ans6_4, A1=>
      nx18619, S0=>nx43185);
   ix31212 : mux21_ni port map ( Y=>nx31211, A0=>max_calc_ans5_4, A1=>
      nx19324, S0=>nx42873);
   ix19325 : mux21 port map ( Y=>nx19324, A0=>nx34896, A1=>nx34903, S0=>
      nx43003);
   ix19385 : xor2 port map ( Y=>nx19384, A0=>nx40661, A1=>
      max_calc_comparator_first_inp1_4);
   ix40698 : xor2 port map ( Y=>nx40697, A0=>
      max_calc_comparator_first_inp2_3, A1=>max_calc_comparator_first_inp1_3
   );
   ix31332 : mux21_ni port map ( Y=>nx31331, A0=>
      max_calc_comparator_first_inp2_3, A1=>nx19498, S0=>nx43397);
   ix19499 : mux21_ni port map ( Y=>nx19498, A0=>nx19494, A1=>nx19406, S0=>
      nx43037);
   ix19407 : mux21_ni port map ( Y=>nx19406, A0=>max_calc_ans2_3, A1=>
      label_2_output_3, S0=>nx43157);
   ix31262 : mux21_ni port map ( Y=>nx31261, A0=>nx19396, A1=>
      max_calc_ans2_3, S0=>nx42997);
   ix19397 : mux21 port map ( Y=>nx19396, A0=>nx40178, A1=>nx40187, S0=>
      nx43021);
   ix19495 : mux21_ni port map ( Y=>nx19494, A0=>max_calc_ans8_3, A1=>
      max_calc_ans7_3, S0=>nx43157);
   ix31322 : mux21_ni port map ( Y=>nx31321, A0=>max_calc_ans7_3, A1=>
      nx19396, S0=>nx43185);
   ix31312 : mux21_ni port map ( Y=>nx31311, A0=>max_calc_ans8_3, A1=>
      nx18620, S0=>nx43287);
   ix19475 : mux21_ni port map ( Y=>nx18620, A0=>
      max_calc_comparator_first_inp2_3, A1=>max_calc_comparator_first_inp1_3, 
      S0=>nx43027);
   ix31302 : mux21_ni port map ( Y=>nx31301, A0=>
      max_calc_comparator_first_inp1_3, A1=>nx19460, S0=>nx43397);
   ix19461 : mux21_ni port map ( Y=>nx19460, A0=>nx19456, A1=>nx19424, S0=>
      nx43037);
   ix19425 : mux21_ni port map ( Y=>nx19424, A0=>max_calc_ans1_3, A1=>
      label_1_output_3, S0=>nx43159);
   ix31272 : mux21_ni port map ( Y=>nx31271, A0=>nx18620, A1=>
      max_calc_ans1_3, S0=>nx42997);
   ix19457 : mux21_ni port map ( Y=>nx19456, A0=>max_calc_ans5_3, A1=>
      max_calc_ans6_3, S0=>nx43159);
   ix31282 : mux21_ni port map ( Y=>nx31281, A0=>max_calc_ans6_3, A1=>
      nx18620, S0=>nx43185);
   ix31292 : mux21_ni port map ( Y=>nx31291, A0=>max_calc_ans5_3, A1=>
      nx19446, S0=>nx42873);
   ix19447 : mux21 port map ( Y=>nx19446, A0=>nx34913, A1=>nx34917, S0=>
      nx43003);
   ix31412 : mux21_ni port map ( Y=>nx31411, A0=>
      max_calc_comparator_first_inp2_2, A1=>nx19620, S0=>nx43397);
   ix19621 : mux21_ni port map ( Y=>nx19620, A0=>nx19616, A1=>nx19528, S0=>
      nx43039);
   ix19529 : mux21_ni port map ( Y=>nx19528, A0=>max_calc_ans2_2, A1=>
      label_2_output_2, S0=>nx43159);
   ix31342 : mux21_ni port map ( Y=>nx31341, A0=>nx19518, A1=>
      max_calc_ans2_2, S0=>nx42997);
   ix19519 : mux21 port map ( Y=>nx19518, A0=>nx40199, A1=>nx40211, S0=>
      nx43021);
   ix19617 : mux21_ni port map ( Y=>nx19616, A0=>max_calc_ans8_2, A1=>
      max_calc_ans7_2, S0=>nx43159);
   ix31402 : mux21_ni port map ( Y=>nx31401, A0=>max_calc_ans7_2, A1=>
      nx19518, S0=>nx43185);
   ix31392 : mux21_ni port map ( Y=>nx31391, A0=>max_calc_ans8_2, A1=>
      nx18621, S0=>nx43287);
   ix19597 : mux21_ni port map ( Y=>nx18621, A0=>
      max_calc_comparator_first_inp2_2, A1=>max_calc_comparator_first_inp1_2, 
      S0=>nx43027);
   ix31382 : mux21_ni port map ( Y=>nx31381, A0=>
      max_calc_comparator_first_inp1_2, A1=>nx19582, S0=>nx43397);
   ix19583 : mux21_ni port map ( Y=>nx19582, A0=>nx19578, A1=>nx19546, S0=>
      nx43039);
   ix19547 : mux21_ni port map ( Y=>nx19546, A0=>max_calc_ans1_2, A1=>
      label_1_output_2, S0=>nx43159);
   ix31352 : mux21_ni port map ( Y=>nx31351, A0=>nx18621, A1=>
      max_calc_ans1_2, S0=>nx42997);
   ix19579 : mux21_ni port map ( Y=>nx19578, A0=>max_calc_ans5_2, A1=>
      max_calc_ans6_2, S0=>nx43159);
   ix31362 : mux21_ni port map ( Y=>nx31361, A0=>max_calc_ans6_2, A1=>
      nx18621, S0=>nx43185);
   ix31372 : mux21_ni port map ( Y=>nx31371, A0=>max_calc_ans5_2, A1=>
      nx19568, S0=>nx42875);
   ix19569 : mux21 port map ( Y=>nx19568, A0=>nx34924, A1=>nx34931, S0=>
      nx43003);
   ix19629 : xor2 port map ( Y=>nx19628, A0=>nx40734, A1=>
      max_calc_comparator_first_inp1_2);
   ix31492 : mux21_ni port map ( Y=>nx31491, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx19742, S0=>nx43399);
   ix19743 : mux21_ni port map ( Y=>nx19742, A0=>nx19738, A1=>nx19650, S0=>
      nx43039);
   ix19651 : mux21_ni port map ( Y=>nx19650, A0=>max_calc_ans2_1, A1=>
      label_2_output_1, S0=>nx43159);
   ix31422 : mux21_ni port map ( Y=>nx31421, A0=>nx19640, A1=>
      max_calc_ans2_1, S0=>nx42997);
   ix19641 : mux21 port map ( Y=>nx19640, A0=>nx40224, A1=>nx40233, S0=>
      nx43021);
   ix19739 : mux21_ni port map ( Y=>nx19738, A0=>max_calc_ans8_1, A1=>
      max_calc_ans7_1, S0=>nx43161);
   ix31482 : mux21_ni port map ( Y=>nx31481, A0=>max_calc_ans7_1, A1=>
      nx19640, S0=>nx43185);
   ix31472 : mux21_ni port map ( Y=>nx31471, A0=>max_calc_ans8_1, A1=>
      nx18622, S0=>nx43289);
   ix19719 : mux21_ni port map ( Y=>nx18622, A0=>
      max_calc_comparator_first_inp2_1, A1=>max_calc_comparator_first_inp1_1, 
      S0=>nx43029);
   ix31462 : mux21_ni port map ( Y=>nx31461, A0=>
      max_calc_comparator_first_inp1_1, A1=>nx19704, S0=>nx43399);
   ix19705 : mux21_ni port map ( Y=>nx19704, A0=>nx19700, A1=>nx19668, S0=>
      nx43039);
   ix19669 : mux21_ni port map ( Y=>nx19668, A0=>max_calc_ans1_1, A1=>
      label_1_output_1, S0=>nx43161);
   ix31432 : mux21_ni port map ( Y=>nx31431, A0=>nx18622, A1=>
      max_calc_ans1_1, S0=>nx42999);
   ix19701 : mux21_ni port map ( Y=>nx19700, A0=>max_calc_ans5_1, A1=>
      max_calc_ans6_1, S0=>nx43161);
   ix31442 : mux21_ni port map ( Y=>nx31441, A0=>max_calc_ans6_1, A1=>
      nx18622, S0=>nx43185);
   ix31452 : mux21_ni port map ( Y=>nx31451, A0=>max_calc_ans5_1, A1=>
      nx19690, S0=>nx42875);
   ix19691 : mux21 port map ( Y=>nx19690, A0=>nx34939, A1=>nx34943, S0=>
      nx43003);
   ix31532 : mux21_ni port map ( Y=>nx31531, A0=>
      max_calc_comparator_first_inp2_0, A1=>nx19800, S0=>nx43399);
   ix19801 : mux21_ni port map ( Y=>nx19800, A0=>nx19796, A1=>nx19772, S0=>
      nx43039);
   ix19773 : mux21_ni port map ( Y=>nx19772, A0=>max_calc_ans2_0, A1=>
      label_2_output_0, S0=>nx43161);
   ix31502 : mux21_ni port map ( Y=>nx31501, A0=>nx19762, A1=>
      max_calc_ans2_0, S0=>nx42999);
   ix19763 : mux21 port map ( Y=>nx19762, A0=>nx40245, A1=>nx40257, S0=>
      nx43023);
   ix19797 : mux21_ni port map ( Y=>nx19796, A0=>max_calc_ans8_0, A1=>
      max_calc_ans7_0, S0=>nx43161);
   ix31522 : mux21_ni port map ( Y=>nx31521, A0=>max_calc_ans7_0, A1=>
      nx19762, S0=>nx43187);
   ix31512 : mux21_ni port map ( Y=>nx31511, A0=>max_calc_ans8_0, A1=>
      nx18213, S0=>nx43289);
   ix20123 : mux21_ni port map ( Y=>nx18213, A0=>
      max_calc_comparator_first_inp2_0, A1=>max_calc_comparator_first_inp1_0, 
      S0=>nx43029);
   ix22882 : mux21_ni port map ( Y=>nx22881, A0=>
      max_calc_comparator_first_inp1_0, A1=>nx6000, S0=>nx43399);
   ix6001 : mux21_ni port map ( Y=>nx6000, A0=>nx5996, A1=>nx2876, S0=>
      nx43039);
   ix2877 : mux21_ni port map ( Y=>nx2876, A0=>max_calc_ans1_0, A1=>
      label_1_output_0, S0=>nx43161);
   ix20832 : mux21_ni port map ( Y=>nx20831, A0=>nx18213, A1=>
      max_calc_ans1_0, S0=>nx42999);
   ix5997 : mux21_ni port map ( Y=>nx5996, A0=>max_calc_ans5_0, A1=>
      max_calc_ans6_0, S0=>nx43161);
   ix20842 : mux21_ni port map ( Y=>nx20841, A0=>max_calc_ans6_0, A1=>
      nx18213, S0=>nx43187);
   ix22872 : mux21_ni port map ( Y=>nx22871, A0=>max_calc_ans5_0, A1=>nx5986, 
      S0=>nx42875);
   ix5987 : mux21 port map ( Y=>nx5986, A0=>nx34950, A1=>nx34957, S0=>
      nx43005);
   ix19751 : xor2 port map ( Y=>nx19750, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx40800);
   ix31652 : mux21_ni port map ( Y=>nx31651, A0=>
      max_calc_comparator_first_inp2_15, A1=>nx20104, S0=>nx43399);
   ix20105 : mux21_ni port map ( Y=>nx20104, A0=>nx20100, A1=>nx19980, S0=>
      nx43039);
   ix19981 : mux21_ni port map ( Y=>nx19980, A0=>max_calc_ans2_15, A1=>
      label_2_output_15, S0=>nx42457);
   ix31552 : mux21_ni port map ( Y=>nx31551, A0=>label_2_output_15, A1=>
      label_2_input_15, S0=>nx42815);
   ix19949 : mux21_ni port map ( Y=>nx19948, A0=>nx19944, A1=>
      label_2_input_state_machine_15, S0=>nx42293);
   ix31542 : mux21_ni port map ( Y=>nx31541, A0=>
      label_2_input_state_machine_15, A1=>data_in(31), S0=>nx42801);
   ix19943 : xnor2 port map ( Y=>nx19942, A0=>nx35419, A1=>label_2_output_15
   );
   ix31562 : mux21_ni port map ( Y=>nx31561, A0=>nx19970, A1=>
      max_calc_ans2_15, S0=>nx42999);
   ix19971 : mux21 port map ( Y=>nx19970, A0=>nx40270, A1=>nx40295, S0=>
      nx43023);
   ix20101 : mux21_ni port map ( Y=>nx20100, A0=>max_calc_ans8_15, A1=>
      max_calc_ans7_15, S0=>nx42457);
   ix31642 : mux21_ni port map ( Y=>nx31641, A0=>max_calc_ans7_15, A1=>
      nx19970, S0=>nx43187);
   ix31632 : mux21_ni port map ( Y=>nx31631, A0=>max_calc_ans8_15, A1=>
      nx18623, S0=>nx43289);
   ix40872 : nor04 port map ( Y=>nx42775, A0=>nx18187, A1=>nx31896, A2=>
      nx43389, A3=>nx42927);
   ix40875 : xor2 port map ( Y=>nx40874, A0=>nx42209, A1=>nx34089);
   ix31792 : mux21_ni port map ( Y=>nx31791, A0=>nx42209, A1=>nx18607, S0=>
      nx43335);
   ix31782 : mux21_ni port map ( Y=>nx31781, A0=>nx42205, A1=>nx18608, S0=>
      nx43335);
   ix40886 : xor2 port map ( Y=>nx40885, A0=>nx42201, A1=>nx34074);
   ix31772 : mux21_ni port map ( Y=>nx31771, A0=>nx42201, A1=>nx18609, S0=>
      nx43335);
   ix31762 : mux21_ni port map ( Y=>nx31761, A0=>nx42197, A1=>nx18610, S0=>
      nx43335);
   ix40896 : xor2 port map ( Y=>nx40895, A0=>nx42193, A1=>nx34059);
   ix31752 : mux21_ni port map ( Y=>nx31751, A0=>nx42193, A1=>nx18611, S0=>
      nx43335);
   ix31742 : mux21_ni port map ( Y=>nx31741, A0=>nx42189, A1=>nx18612, S0=>
      nx43337);
   ix40907 : xor2 port map ( Y=>nx40906, A0=>nx42185, A1=>nx34044);
   ix31732 : mux21_ni port map ( Y=>nx31731, A0=>nx42185, A1=>nx18613, S0=>
      nx43337);
   ix31722 : mux21_ni port map ( Y=>nx31721, A0=>nx42181, A1=>nx18615, S0=>
      nx43337);
   ix40917 : xor2 port map ( Y=>nx40916, A0=>nx42177, A1=>nx34029);
   ix31712 : mux21_ni port map ( Y=>nx31711, A0=>nx42177, A1=>nx18617, S0=>
      nx43337);
   ix31702 : mux21_ni port map ( Y=>nx31701, A0=>nx42173, A1=>nx18619, S0=>
      nx43337);
   ix40928 : xor2 port map ( Y=>nx40927, A0=>nx42169, A1=>nx34014);
   ix31692 : mux21_ni port map ( Y=>nx31691, A0=>nx42169, A1=>nx18620, S0=>
      nx43337);
   ix31682 : mux21_ni port map ( Y=>nx31681, A0=>nx42165, A1=>nx18621, S0=>
      nx43337);
   ix40938 : xor2 port map ( Y=>nx40937, A0=>nx42161, A1=>nx33999);
   ix31672 : mux21_ni port map ( Y=>nx31671, A0=>nx42161, A1=>nx18622, S0=>
      nx43339);
   ix31662 : mux21_ni port map ( Y=>nx31661, A0=>nx41531, A1=>nx18213, S0=>
      nx43339);
   ix40951 : xor2 port map ( Y=>nx40950, A0=>nx42217, A1=>nx34987);
   ix40955 : xor2 port map ( Y=>nx40954, A0=>nx42209, A1=>nx34754);
   ix40960 : xor2 port map ( Y=>nx40959, A0=>nx42201, A1=>nx34739);
   ix40964 : xor2 port map ( Y=>nx40963, A0=>nx42193, A1=>nx34724);
   ix40969 : xor2 port map ( Y=>nx40968, A0=>nx42185, A1=>nx34709);
   ix40973 : xor2 port map ( Y=>nx40972, A0=>nx42177, A1=>nx34694);
   ix40978 : xor2 port map ( Y=>nx40977, A0=>nx42169, A1=>nx34679);
   ix40982 : xor2 port map ( Y=>nx40981, A0=>nx42161, A1=>nx34664);
   ix40986 : or04 port map ( Y=>nx40985, A0=>nx43389, A1=>nx42927, A2=>
      nx33436, A3=>nx43453);
   ix20063 : mux21_ni port map ( Y=>nx20062, A0=>max_calc_ans5_15, A1=>
      max_calc_ans6_15, S0=>nx42457);
   ix31602 : mux21_ni port map ( Y=>nx31601, A0=>max_calc_ans6_15, A1=>
      nx18623, S0=>nx43187);
   ix31612 : mux21_ni port map ( Y=>nx31611, A0=>max_calc_ans5_15, A1=>
      nx20052, S0=>nx42875);
   ix20053 : mux21 port map ( Y=>nx20052, A0=>nx34965, A1=>nx34971, S0=>
      nx43005);
   ix41001 : xor2 port map ( Y=>nx41000, A0=>nx42209, A1=>nx39051);
   ix41006 : xor2 port map ( Y=>nx41005, A0=>nx42201, A1=>nx39036);
   ix41010 : xor2 port map ( Y=>nx41009, A0=>nx42193, A1=>nx39021);
   ix41015 : xor2 port map ( Y=>nx41014, A0=>nx42185, A1=>nx39006);
   ix41019 : xor2 port map ( Y=>nx41018, A0=>nx42177, A1=>nx38991);
   ix41024 : xor2 port map ( Y=>nx41023, A0=>nx42169, A1=>nx38976);
   ix41028 : xor2 port map ( Y=>nx41027, A0=>nx42161, A1=>nx38961);
   ix41039 : xor2 port map ( Y=>nx41038, A0=>nx42161, A1=>nx37445);
   ix41043 : xor2 port map ( Y=>nx41042, A0=>nx42169, A1=>nx37460);
   ix41049 : xor2 port map ( Y=>nx41048, A0=>nx42177, A1=>nx37475);
   ix41053 : xor2 port map ( Y=>nx41052, A0=>nx42185, A1=>nx37490);
   ix41059 : xor2 port map ( Y=>nx41058, A0=>nx42193, A1=>nx37505);
   ix41063 : xor2 port map ( Y=>nx41062, A0=>nx42201, A1=>nx37520);
   ix41069 : xor2 port map ( Y=>nx41068, A0=>nx42209, A1=>nx37535);
   ix41073 : xor2 port map ( Y=>nx41072, A0=>nx42217, A1=>nx37756);
   ix41081 : xor2 port map ( Y=>nx41080, A0=>nx42217, A1=>nx40312);
   ix41085 : xor2 port map ( Y=>nx41084, A0=>nx42209, A1=>nx36262);
   ix41090 : xor2 port map ( Y=>nx41089, A0=>nx42201, A1=>nx36247);
   ix41094 : xor2 port map ( Y=>nx41093, A0=>nx42193, A1=>nx36232);
   ix41099 : xor2 port map ( Y=>nx41098, A0=>nx42185, A1=>nx36217);
   ix41103 : xor2 port map ( Y=>nx41102, A0=>nx42177, A1=>nx36202);
   ix41108 : xor2 port map ( Y=>nx41107, A0=>nx42169, A1=>nx36187);
   ix41112 : xor2 port map ( Y=>nx41111, A0=>nx42161, A1=>nx36172);
   ix41123 : xor2 port map ( Y=>nx41122, A0=>nx42161, A1=>nx35534);
   ix41127 : xor2 port map ( Y=>nx41126, A0=>nx42169, A1=>nx35549);
   ix41133 : xor2 port map ( Y=>nx41132, A0=>nx42177, A1=>nx35564);
   ix41137 : xor2 port map ( Y=>nx41136, A0=>nx42185, A1=>nx35579);
   ix41143 : xor2 port map ( Y=>nx41142, A0=>nx42193, A1=>nx35594);
   ix41147 : xor2 port map ( Y=>nx41146, A0=>nx42201, A1=>nx35609);
   ix41153 : xor2 port map ( Y=>nx41152, A0=>nx42209, A1=>nx35624);
   ix41157 : xor2 port map ( Y=>nx41156, A0=>nx42217, A1=>nx40857);
   ix41162 : xor2 port map ( Y=>nx41161, A0=>nx42219, A1=>nx33421);
   ix41166 : xor2 port map ( Y=>nx41165, A0=>nx42211, A1=>nx33415);
   ix41171 : xor2 port map ( Y=>nx41170, A0=>nx42203, A1=>nx33400);
   ix41175 : xor2 port map ( Y=>nx41174, A0=>nx42195, A1=>nx33385);
   ix41180 : xor2 port map ( Y=>nx41179, A0=>nx42187, A1=>nx33370);
   ix41184 : xor2 port map ( Y=>nx41183, A0=>nx42179, A1=>nx33355);
   ix41189 : xor2 port map ( Y=>nx41188, A0=>nx42171, A1=>nx33340);
   ix41193 : xor2 port map ( Y=>nx41192, A0=>nx42163, A1=>nx33325);
   ix41199 : xor2 port map ( Y=>nx41198, A0=>nx42219, A1=>nx40287);
   ix41203 : xor2 port map ( Y=>nx41202, A0=>nx42211, A1=>nx38414);
   ix41208 : xor2 port map ( Y=>nx41207, A0=>nx42203, A1=>nx38399);
   ix41212 : xor2 port map ( Y=>nx41211, A0=>nx42195, A1=>nx38384);
   ix41217 : xor2 port map ( Y=>nx41216, A0=>nx42187, A1=>nx38369);
   ix41221 : xor2 port map ( Y=>nx41220, A0=>nx42179, A1=>nx38354);
   ix41226 : xor2 port map ( Y=>nx41225, A0=>nx42171, A1=>nx38339);
   ix41230 : xor2 port map ( Y=>nx41229, A0=>nx42163, A1=>nx38324);
   ix41237 : xor2 port map ( Y=>nx41236, A0=>nx42219, A1=>nx37776);
   ix41241 : xor2 port map ( Y=>nx41240, A0=>nx42211, A1=>nx36899);
   ix41246 : xor2 port map ( Y=>nx41245, A0=>nx42203, A1=>nx36884);
   ix41250 : xor2 port map ( Y=>nx41249, A0=>nx42195, A1=>nx36869);
   ix41255 : xor2 port map ( Y=>nx41254, A0=>nx42187, A1=>nx36854);
   ix41259 : xor2 port map ( Y=>nx41258, A0=>nx42179, A1=>nx36839);
   ix41264 : xor2 port map ( Y=>nx41263, A0=>nx42171, A1=>nx36824);
   ix41268 : xor2 port map ( Y=>nx41267, A0=>nx42163, A1=>nx36809);
   ix41274 : xor2 port map ( Y=>nx41273, A0=>nx42219, A1=>nx39906);
   ix41278 : xor2 port map ( Y=>nx41277, A0=>nx42211, A1=>nx39685);
   ix41283 : xor2 port map ( Y=>nx41282, A0=>nx42203, A1=>nx39670);
   ix41287 : xor2 port map ( Y=>nx41286, A0=>nx42195, A1=>nx39655);
   ix41292 : xor2 port map ( Y=>nx41291, A0=>nx42187, A1=>nx39640);
   ix41296 : xor2 port map ( Y=>nx41295, A0=>nx42179, A1=>nx39625);
   ix41301 : xor2 port map ( Y=>nx41300, A0=>nx42171, A1=>nx39610);
   ix41305 : xor2 port map ( Y=>nx41304, A0=>nx42163, A1=>nx39595);
   ix41314 : and02 port map ( Y=>nx41313, A0=>nx42247, A1=>nx42927);
   ix41322 : nor02ii port map ( Y=>nx41321, A0=>nx41325, A1=>nx32709);
   ix1613 : nor02ii port map ( Y=>nx1612, A0=>nx41354, A1=>nx42863);
   ix21063 : and04 port map ( Y=>nx21062, A0=>sub_state_2, A1=>nx42863, A2=>
      nx42869, A3=>nx42881);
   ix21047 : ao21 port map ( Y=>nx21046, A0=>nx42869, A1=>nx42881, B0=>
      nx42257);
   ix42846 : inv02 port map ( Y=>nx42847, A=>nx42249);
   ix42848 : inv02 port map ( Y=>nx42849, A=>nx42249);
   ix42850 : inv02 port map ( Y=>nx42851, A=>nx42249);
   ix42852 : inv02 port map ( Y=>nx42853, A=>nx42249);
   ix42854 : inv02 port map ( Y=>nx42855, A=>nx42277);
   ix42856 : inv02 port map ( Y=>nx42857, A=>nx42277);
   ix42858 : inv02 port map ( Y=>nx42859, A=>nx42277);
   ix42860 : inv02 port map ( Y=>nx42861, A=>nx42893);
   ix42862 : inv02 port map ( Y=>nx42863, A=>nx42893);
   ix42864 : inv02 port map ( Y=>nx42865, A=>nx41360);
   ix42866 : inv02 port map ( Y=>nx42867, A=>nx42273);
   ix42868 : inv02 port map ( Y=>nx42869, A=>nx42273);
   ix42870 : inv02 port map ( Y=>nx42871, A=>nx42527);
   ix42872 : inv02 port map ( Y=>nx42873, A=>nx42527);
   ix42874 : inv02 port map ( Y=>nx42875, A=>nx42527);
   ix42876 : inv02 port map ( Y=>nx42877, A=>state_2);
   ix42878 : inv02 port map ( Y=>nx42879, A=>state_2);
   ix42880 : inv02 port map ( Y=>nx42881, A=>nx41381);
   ix42882 : inv02 port map ( Y=>nx42883, A=>nx41383);
   ix42884 : inv02 port map ( Y=>nx42885, A=>nx41383);
   ix42886 : inv02 port map ( Y=>nx42887, A=>nx41405);
   ix42888 : inv02 port map ( Y=>nx42889, A=>nx41405);
   ix42890 : inv02 port map ( Y=>nx42891, A=>sub_state_0);
   ix42892 : inv02 port map ( Y=>nx42893, A=>sub_state_0);
   ix42894 : inv01 port map ( Y=>nx42895, A=>nx31985);
   ix42896 : inv02 port map ( Y=>nx42897, A=>nx42895);
   ix42898 : inv02 port map ( Y=>nx42899, A=>nx42895);
   ix42900 : inv02 port map ( Y=>nx42901, A=>nx42895);
   ix42902 : inv02 port map ( Y=>nx42903, A=>nx42895);
   ix42904 : inv01 port map ( Y=>nx42905, A=>nx32101);
   ix42906 : inv02 port map ( Y=>nx42907, A=>nx42905);
   ix42908 : inv02 port map ( Y=>nx42909, A=>nx42905);
   ix42910 : inv02 port map ( Y=>nx42911, A=>nx42905);
   ix42912 : inv01 port map ( Y=>nx42913, A=>nx32142);
   ix42914 : inv02 port map ( Y=>nx42915, A=>nx42913);
   ix42916 : inv02 port map ( Y=>nx42917, A=>nx42913);
   ix42918 : inv02 port map ( Y=>nx42919, A=>nx42913);
   ix42920 : buf02 port map ( Y=>nx42921, A=>nx32886);
   ix42922 : buf02 port map ( Y=>nx42923, A=>nx32886);
   ix42924 : inv02 port map ( Y=>nx42925, A=>nx41371);
   ix42926 : inv02 port map ( Y=>nx42927, A=>nx41371);
   ix42928 : buf02 port map ( Y=>nx42929, A=>nx33610);
   ix42930 : buf02 port map ( Y=>nx42931, A=>nx33610);
   ix42932 : buf02 port map ( Y=>nx42933, A=>nx34275);
   ix42934 : buf02 port map ( Y=>nx42935, A=>nx34275);
   ix42936 : buf02 port map ( Y=>nx42937, A=>nx35145);
   ix42938 : buf02 port map ( Y=>nx42939, A=>nx35145);
   ix42940 : buf02 port map ( Y=>nx42941, A=>nx35783);
   ix42942 : buf02 port map ( Y=>nx42943, A=>nx35783);
   ix42944 : buf02 port map ( Y=>nx42945, A=>nx36420);
   ix42946 : buf02 port map ( Y=>nx42947, A=>nx36420);
   ix42948 : buf02 port map ( Y=>nx42949, A=>nx37056);
   ix42950 : buf02 port map ( Y=>nx42951, A=>nx37056);
   ix42952 : buf02 port map ( Y=>nx42953, A=>nx37935);
   ix42954 : buf02 port map ( Y=>nx42955, A=>nx37935);
   ix42956 : buf02 port map ( Y=>nx42957, A=>nx38572);
   ix42958 : buf02 port map ( Y=>nx42959, A=>nx38572);
   ix42960 : buf02 port map ( Y=>nx42961, A=>nx39206);
   ix42962 : buf02 port map ( Y=>nx42963, A=>nx39206);
   ix42964 : inv02 port map ( Y=>nx42965, A=>nx294);
   ix42966 : inv02 port map ( Y=>nx42967, A=>nx294);
   ix42968 : inv02 port map ( Y=>nx42969, A=>nx294);
   ix42970 : inv02 port map ( Y=>nx42971, A=>nx41523);
   ix42972 : inv02 port map ( Y=>nx42973, A=>nx41523);
   ix42974 : inv02 port map ( Y=>nx42975, A=>nx41577);
   ix42976 : inv02 port map ( Y=>nx42977, A=>nx41577);
   ix42978 : inv02 port map ( Y=>nx42979, A=>nx41577);
   ix42980 : inv01 port map ( Y=>nx42981, A=>nx41733);
   ix42982 : inv02 port map ( Y=>nx42983, A=>nx42981);
   ix42984 : inv02 port map ( Y=>nx42985, A=>nx42981);
   ix42986 : inv02 port map ( Y=>nx42987, A=>nx42981);
   ix42988 : inv01 port map ( Y=>nx42989, A=>nx41821);
   ix42990 : inv02 port map ( Y=>nx42991, A=>nx42989);
   ix42992 : inv02 port map ( Y=>nx42993, A=>nx42989);
   ix42994 : inv02 port map ( Y=>nx42995, A=>nx42989);
   ix42996 : inv02 port map ( Y=>nx42997, A=>nx42989);
   ix42998 : inv02 port map ( Y=>nx42999, A=>nx42989);
   ix43000 : inv02 port map ( Y=>nx43001, A=>nx5978);
   ix43002 : inv02 port map ( Y=>nx43003, A=>nx5978);
   ix43004 : inv02 port map ( Y=>nx43005, A=>nx5978);
   ix43006 : inv02 port map ( Y=>nx43007, A=>nx11786);
   ix43008 : inv02 port map ( Y=>nx43009, A=>nx11786);
   ix43010 : inv02 port map ( Y=>nx43011, A=>nx11786);
   ix43012 : inv02 port map ( Y=>nx43013, A=>nx16276);
   ix43014 : inv02 port map ( Y=>nx43015, A=>nx16276);
   ix43016 : inv02 port map ( Y=>nx43017, A=>nx16276);
   ix43018 : inv02 port map ( Y=>nx43019, A=>nx17604);
   ix43020 : inv02 port map ( Y=>nx43021, A=>nx17604);
   ix43022 : inv02 port map ( Y=>nx43023, A=>nx17604);
   ix43024 : inv02 port map ( Y=>nx43025, A=>nx18605);
   ix43026 : inv02 port map ( Y=>nx43027, A=>nx18605);
   ix43028 : inv02 port map ( Y=>nx43029, A=>nx18605);
   ix43030 : inv02 port map ( Y=>nx43031, A=>nx43389);
   ix43032 : inv02 port map ( Y=>nx43033, A=>nx42805);
   ix43034 : inv02 port map ( Y=>nx43035, A=>nx42805);
   ix43036 : inv02 port map ( Y=>nx43037, A=>nx42805);
   ix43038 : inv02 port map ( Y=>nx43039, A=>nx42805);
   ix43040 : inv02 port map ( Y=>nx43041, A=>sub_state_2);
   ix43042 : inv02 port map ( Y=>nx43043, A=>sub_state_2);
   ix43044 : inv02 port map ( Y=>nx43045, A=>sub_state_2);
   ix43046 : inv01 port map ( Y=>nx43047, A=>nx42263);
   ix43048 : inv02 port map ( Y=>nx43049, A=>nx43047);
   ix43050 : inv02 port map ( Y=>nx43051, A=>nx43047);
   ix43052 : inv02 port map ( Y=>nx43053, A=>nx43047);
   ix43054 : inv02 port map ( Y=>nx43055, A=>nx43445);
   ix43056 : inv02 port map ( Y=>nx43057, A=>nx43445);
   ix43058 : inv02 port map ( Y=>nx43059, A=>nx43445);
   ix43060 : inv02 port map ( Y=>nx43061, A=>nx43447);
   ix43062 : inv02 port map ( Y=>nx43063, A=>nx43447);
   ix43064 : inv02 port map ( Y=>nx43065, A=>nx43447);
   ix43066 : inv02 port map ( Y=>nx43067, A=>nx43447);
   ix43068 : inv02 port map ( Y=>nx43069, A=>nx43447);
   ix43070 : inv02 port map ( Y=>nx43071, A=>nx43447);
   ix43072 : inv02 port map ( Y=>nx43073, A=>nx43447);
   ix43074 : inv02 port map ( Y=>nx43075, A=>nx43449);
   ix43076 : inv02 port map ( Y=>nx43077, A=>nx43449);
   ix43078 : inv02 port map ( Y=>nx43079, A=>nx43449);
   ix43080 : inv02 port map ( Y=>nx43081, A=>nx43449);
   ix43082 : inv02 port map ( Y=>nx43083, A=>nx43449);
   ix43084 : inv02 port map ( Y=>nx43085, A=>nx43449);
   ix43086 : inv02 port map ( Y=>nx43087, A=>nx43449);
   ix43088 : inv02 port map ( Y=>nx43089, A=>nx43451);
   ix43090 : inv02 port map ( Y=>nx43091, A=>nx43451);
   ix43092 : inv02 port map ( Y=>nx43093, A=>nx43451);
   ix43094 : inv02 port map ( Y=>nx43095, A=>nx43451);
   ix43096 : inv04 port map ( Y=>nx43097, A=>alu_sel);
   ix43098 : inv04 port map ( Y=>nx43099, A=>alu_sel);
   ix43100 : inv04 port map ( Y=>nx43101, A=>alu_sel);
   ix43102 : inv02 port map ( Y=>nx43103, A=>nx68);
   ix43104 : inv01 port map ( Y=>nx43105, A=>nx42303);
   ix43106 : inv02 port map ( Y=>nx43107, A=>nx43105);
   ix43108 : inv02 port map ( Y=>nx43109, A=>nx43105);
   ix43110 : inv02 port map ( Y=>nx43111, A=>nx43105);
   ix43112 : inv02 port map ( Y=>nx43113, A=>nx42313);
   ix43114 : inv02 port map ( Y=>nx43115, A=>nx42313);
   ix43116 : inv02 port map ( Y=>nx43117, A=>nx32131);
   ix43118 : inv02 port map ( Y=>nx43119, A=>nx32131);
   ix43120 : inv02 port map ( Y=>nx43121, A=>nx32131);
   ix43122 : inv02 port map ( Y=>nx43123, A=>nx43463);
   ix43124 : inv02 port map ( Y=>nx43125, A=>nx43463);
   ix43126 : inv02 port map ( Y=>nx43127, A=>nx43465);
   ix43128 : inv02 port map ( Y=>nx43129, A=>nx43465);
   ix43130 : inv02 port map ( Y=>nx43131, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix43132 : inv02 port map ( Y=>nx43133, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix43134 : inv02 port map ( Y=>nx43135, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix43136 : inv02 port map ( Y=>nx43137, A=>nx43453);
   ix43138 : inv02 port map ( Y=>nx43139, A=>nx43453);
   ix43140 : inv02 port map ( Y=>nx43141, A=>nx43455);
   ix43142 : inv02 port map ( Y=>nx43143, A=>nx43455);
   ix43144 : inv02 port map ( Y=>nx43145, A=>nx43455);
   ix43146 : inv02 port map ( Y=>nx43147, A=>nx43455);
   ix43148 : inv02 port map ( Y=>nx43149, A=>nx43455);
   ix43150 : inv02 port map ( Y=>nx43151, A=>nx43455);
   ix43152 : inv02 port map ( Y=>nx43153, A=>nx43455);
   ix43154 : inv02 port map ( Y=>nx43155, A=>nx43457);
   ix43156 : inv02 port map ( Y=>nx43157, A=>nx43457);
   ix43158 : inv02 port map ( Y=>nx43159, A=>nx43457);
   ix43160 : inv02 port map ( Y=>nx43161, A=>nx43457);
   ix43162 : inv02 port map ( Y=>nx43163, A=>nx43471);
   ix43164 : inv02 port map ( Y=>nx43165, A=>nx43471);
   ix43166 : inv02 port map ( Y=>nx43167, A=>nx43473);
   ix43168 : inv02 port map ( Y=>nx43169, A=>nx43473);
   ix43170 : inv02 port map ( Y=>nx43171, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix43172 : inv02 port map ( Y=>nx43173, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix43174 : inv02 port map ( Y=>nx43175, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix43176 : inv01 port map ( Y=>nx43177, A=>nx42485);
   ix43178 : inv02 port map ( Y=>nx43179, A=>nx43177);
   ix43180 : inv02 port map ( Y=>nx43181, A=>nx43177);
   ix43182 : inv02 port map ( Y=>nx43183, A=>nx43177);
   ix43184 : inv02 port map ( Y=>nx43185, A=>nx43177);
   ix43186 : inv02 port map ( Y=>nx43187, A=>nx43177);
   ix43188 : inv02 port map ( Y=>nx43189, A=>nx43467);
   ix43190 : inv02 port map ( Y=>nx43191, A=>nx43467);
   ix43192 : inv02 port map ( Y=>nx43193, A=>nx43469);
   ix43194 : inv02 port map ( Y=>nx43195, A=>nx43469);
   ix43196 : inv02 port map ( Y=>nx43197, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix43198 : inv02 port map ( Y=>nx43199, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix43200 : inv02 port map ( Y=>nx43201, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix43202 : inv02 port map ( Y=>nx43203, A=>nx2862);
   ix43204 : inv02 port map ( Y=>nx43205, A=>nx43459);
   ix43206 : inv02 port map ( Y=>nx43207, A=>nx43459);
   ix43208 : inv02 port map ( Y=>nx43209, A=>nx43461);
   ix43210 : inv02 port map ( Y=>nx43211, A=>nx43461);
   ix43212 : inv02 port map ( Y=>nx43213, A=>nx43461);
   ix43214 : inv02 port map ( Y=>nx43215, A=>nx43461);
   ix43216 : inv02 port map ( Y=>nx43217, A=>nx43461);
   ix43218 : inv02 port map ( Y=>nx43219, A=>nx43461);
   ix43220 : inv02 port map ( Y=>nx43221, A=>nx43475);
   ix43222 : inv02 port map ( Y=>nx43223, A=>nx43475);
   ix43224 : inv02 port map ( Y=>nx43225, A=>nx43477);
   ix43226 : inv02 port map ( Y=>nx43227, A=>nx43477);
   ix43228 : inv02 port map ( Y=>nx43229, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix43230 : inv02 port map ( Y=>nx43231, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix43232 : inv02 port map ( Y=>nx43233, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix43234 : inv02 port map ( Y=>nx43235, A=>nx43479);
   ix43236 : inv02 port map ( Y=>nx43237, A=>nx43479);
   ix43238 : inv02 port map ( Y=>nx43239, A=>nx43481);
   ix43240 : inv02 port map ( Y=>nx43241, A=>nx43481);
   ix43242 : inv02 port map ( Y=>nx43243, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix43244 : inv02 port map ( Y=>nx43245, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix43246 : inv02 port map ( Y=>nx43247, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix43248 : inv02 port map ( Y=>nx43249, A=>nx43483);
   ix43250 : inv02 port map ( Y=>nx43251, A=>nx43483);
   ix43252 : inv02 port map ( Y=>nx43253, A=>nx43485);
   ix43254 : inv02 port map ( Y=>nx43255, A=>nx43485);
   ix43256 : inv02 port map ( Y=>nx43257, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix43258 : inv02 port map ( Y=>nx43259, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix43260 : inv02 port map ( Y=>nx43261, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix43262 : inv02 port map ( Y=>nx43263, A=>nx36903);
   ix43264 : inv02 port map ( Y=>nx43265, A=>nx36903);
   ix43266 : inv02 port map ( Y=>nx43267, A=>nx36903);
   ix43268 : inv02 port map ( Y=>nx43269, A=>nx43487);
   ix43270 : inv02 port map ( Y=>nx43271, A=>nx43487);
   ix43272 : inv02 port map ( Y=>nx43273, A=>nx43489);
   ix43274 : inv02 port map ( Y=>nx43275, A=>nx43489);
   ix43276 : inv02 port map ( Y=>nx43277, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix43278 : inv02 port map ( Y=>nx43279, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix43280 : inv02 port map ( Y=>nx43281, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix43282 : inv01 port map ( Y=>nx43283, A=>nx42689);
   ix43284 : inv02 port map ( Y=>nx43285, A=>nx43283);
   ix43286 : inv02 port map ( Y=>nx43287, A=>nx43283);
   ix43288 : inv02 port map ( Y=>nx43289, A=>nx43283);
   ix43290 : inv02 port map ( Y=>nx43291, A=>nx43491);
   ix43292 : inv02 port map ( Y=>nx43293, A=>nx43491);
   ix43294 : inv02 port map ( Y=>nx43295, A=>nx43493);
   ix43296 : inv02 port map ( Y=>nx43297, A=>nx43493);
   ix43298 : inv02 port map ( Y=>nx43299, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix43300 : inv02 port map ( Y=>nx43301, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix43302 : inv02 port map ( Y=>nx43303, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix43304 : inv02 port map ( Y=>nx43305, A=>nx43495);
   ix43306 : inv02 port map ( Y=>nx43307, A=>nx43495);
   ix43308 : inv02 port map ( Y=>nx43309, A=>nx43497);
   ix43310 : inv02 port map ( Y=>nx43311, A=>nx43497);
   ix43312 : inv02 port map ( Y=>nx43313, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix43314 : inv02 port map ( Y=>nx43315, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix43316 : inv02 port map ( Y=>nx43317, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix43318 : inv02 port map ( Y=>nx43319, A=>nx43499);
   ix43320 : inv02 port map ( Y=>nx43321, A=>nx43499);
   ix43322 : inv02 port map ( Y=>nx43323, A=>nx43501);
   ix43324 : inv02 port map ( Y=>nx43325, A=>nx43501);
   ix43326 : inv02 port map ( Y=>nx43327, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix43328 : inv02 port map ( Y=>nx43329, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix43330 : inv02 port map ( Y=>nx43331, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix43332 : inv01 port map ( Y=>nx43333, A=>nx42775);
   ix43334 : inv02 port map ( Y=>nx43335, A=>nx43333);
   ix43336 : inv02 port map ( Y=>nx43337, A=>nx43333);
   ix43338 : inv02 port map ( Y=>nx43339, A=>nx43333);
   ix43340 : inv02 port map ( Y=>nx43341, A=>nx36903);
   ix43342 : inv02 port map ( Y=>nx43343, A=>nx36903);
   ix43344 : inv02 port map ( Y=>nx43345, A=>nx36903);
   ix43346 : inv02 port map ( Y=>nx43347, A=>nx36903);
   ix43348 : inv02 port map ( Y=>nx43349, A=>nx43503);
   ix43350 : inv02 port map ( Y=>nx43351, A=>nx43503);
   ix43352 : inv02 port map ( Y=>nx43353, A=>nx43503);
   ix43354 : inv02 port map ( Y=>nx43355, A=>nx43503);
   ix43356 : inv02 port map ( Y=>nx43357, A=>nx43505);
   ix43358 : inv02 port map ( Y=>nx43359, A=>nx43505);
   ix43360 : inv02 port map ( Y=>nx43361, A=>nx43505);
   ix43362 : inv02 port map ( Y=>nx43363, A=>nx43505);
   ix43364 : inv02 port map ( Y=>nx43365, A=>nx43505);
   ix43366 : inv02 port map ( Y=>nx43367, A=>nx43505);
   ix43368 : inv02 port map ( Y=>nx43369, A=>nx43505);
   ix43370 : inv02 port map ( Y=>nx43371, A=>nx43507);
   ix43372 : inv02 port map ( Y=>nx43373, A=>nx43507);
   ix43374 : inv02 port map ( Y=>nx43375, A=>nx43507);
   ix43376 : inv02 port map ( Y=>nx43377, A=>nx43507);
   ix43378 : inv02 port map ( Y=>nx43379, A=>nx43507);
   ix43380 : inv02 port map ( Y=>nx43381, A=>nx43507);
   ix43382 : inv02 port map ( Y=>nx43383, A=>nx43507);
   ix43384 : inv02 port map ( Y=>nx43385, A=>nx43509);
   ix43386 : inv02 port map ( Y=>nx43387, A=>nx43509);
   ix43388 : inv02 port map ( Y=>nx43389, A=>nx42227);
   ix43390 : inv02 port map ( Y=>nx43391, A=>nx34993);
   ix43392 : inv02 port map ( Y=>nx43393, A=>nx34993);
   ix43394 : inv02 port map ( Y=>nx43395, A=>nx34993);
   ix43396 : inv02 port map ( Y=>nx43397, A=>nx34993);
   ix43398 : inv02 port map ( Y=>nx43399, A=>nx34993);
   ix43400 : inv02 port map ( Y=>nx43401, A=>nx43511);
   ix43402 : inv02 port map ( Y=>nx43403, A=>nx43511);
   ix43404 : inv02 port map ( Y=>nx43405, A=>nx43511);
   ix43406 : inv02 port map ( Y=>nx43407, A=>nx43511);
   ix43408 : inv02 port map ( Y=>nx43409, A=>nx43513);
   ix43410 : inv02 port map ( Y=>nx43411, A=>nx43513);
   ix43412 : inv02 port map ( Y=>nx43413, A=>nx43513);
   ix43414 : inv02 port map ( Y=>nx43415, A=>nx43513);
   ix43416 : inv02 port map ( Y=>nx43417, A=>nx43513);
   ix43418 : inv02 port map ( Y=>nx43419, A=>nx43513);
   ix43420 : inv02 port map ( Y=>nx43421, A=>nx43513);
   ix43422 : inv02 port map ( Y=>nx43423, A=>nx43515);
   ix43424 : inv02 port map ( Y=>nx43425, A=>nx43515);
   ix43426 : inv02 port map ( Y=>nx43427, A=>nx43515);
   ix43428 : inv02 port map ( Y=>nx43429, A=>nx43515);
   ix43430 : inv02 port map ( Y=>nx43431, A=>nx43515);
   ix43432 : inv02 port map ( Y=>nx43433, A=>nx43515);
   ix43434 : inv02 port map ( Y=>nx43435, A=>nx43515);
   ix43436 : inv02 port map ( Y=>nx43437, A=>nx43517);
   ix43438 : inv02 port map ( Y=>nx43439, A=>nx43517);
   ix43444 : inv02 port map ( Y=>nx43445, A=>nx42285);
   ix43446 : inv02 port map ( Y=>nx43447, A=>nx42285);
   ix43448 : inv02 port map ( Y=>nx43449, A=>nx42285);
   ix43450 : inv02 port map ( Y=>nx43451, A=>nx42285);
   ix43452 : inv02 port map ( Y=>nx43453, A=>nx42453);
   ix43454 : inv02 port map ( Y=>nx43455, A=>nx42453);
   ix43456 : inv02 port map ( Y=>nx43457, A=>nx42453);
   ix43458 : inv02 port map ( Y=>nx43459, A=>nx34993);
   ix43460 : inv02 port map ( Y=>nx43461, A=>nx34993);
   ix43462 : inv02 port map ( Y=>nx43463, A=>nx42373);
   ix43464 : inv02 port map ( Y=>nx43465, A=>nx42373);
   ix43466 : inv02 port map ( Y=>nx43467, A=>nx42497);
   ix43468 : inv02 port map ( Y=>nx43469, A=>nx42497);
   ix43470 : inv02 port map ( Y=>nx43471, A=>nx42459);
   ix43472 : inv02 port map ( Y=>nx43473, A=>nx42459);
   ix43474 : inv02 port map ( Y=>nx43475, A=>nx42551);
   ix43476 : inv02 port map ( Y=>nx43477, A=>nx42551);
   ix43478 : inv02 port map ( Y=>nx43479, A=>nx42577);
   ix43480 : inv02 port map ( Y=>nx43481, A=>nx42577);
   ix43482 : inv02 port map ( Y=>nx43483, A=>nx42603);
   ix43484 : inv02 port map ( Y=>nx43485, A=>nx42603);
   ix43486 : inv02 port map ( Y=>nx43487, A=>nx42651);
   ix43488 : inv02 port map ( Y=>nx43489, A=>nx42651);
   ix43490 : inv02 port map ( Y=>nx43491, A=>nx42697);
   ix43492 : inv02 port map ( Y=>nx43493, A=>nx42697);
   ix43494 : inv02 port map ( Y=>nx43495, A=>nx42723);
   ix43496 : inv02 port map ( Y=>nx43497, A=>nx42723);
   ix43498 : inv02 port map ( Y=>nx43499, A=>nx42749);
   ix43500 : inv02 port map ( Y=>nx43501, A=>nx42749);
   ix43502 : inv02 port map ( Y=>nx43503, A=>nx42795);
   ix43504 : inv02 port map ( Y=>nx43505, A=>nx42795);
   ix43506 : inv02 port map ( Y=>nx43507, A=>nx42795);
   ix43508 : inv02 port map ( Y=>nx43509, A=>nx42795);
   ix43510 : inv02 port map ( Y=>nx43511, A=>nx42809);
   ix43512 : inv02 port map ( Y=>nx43513, A=>nx42809);
   ix43514 : inv02 port map ( Y=>nx43515, A=>nx42809);
   ix43516 : inv02 port map ( Y=>nx43517, A=>nx42809);
   ix43518 : inv02 port map ( Y=>nx43519, A=>enable_decoder_dst_booth);
   ix43520 : inv02 port map ( Y=>nx43521, A=>nx33312);
end a_FC_controller ;


