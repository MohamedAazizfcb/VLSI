//
// Verilog description for cell IOCHIP, 
// Wed Apr 24 13:15:28 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module IOCHIP ( OuterRead, OuterWrite, ActivateOuterAddress, INCEnable, PDone, 
                OuterAddress, ResultIn, CLK, LP, INTR, CNNIMGLOAD, Rst, 
                EnableReadingFromCPU, DecompressionDone, DecompressionDone1, 
                DecompressionDone2, readenable, DataBus, Address, 
                DecompressedData, DecompressedData1, DecompressedData2, 
                EnableReadingFromCPU1, EnableReadingFromCPU2, loadingimg, 
                loadingCNN, PClk, DataFromRam, Result, Done, ProcessEnable ) ;

    input OuterRead ;
    input OuterWrite ;
    input ActivateOuterAddress ;
    input INCEnable ;
    input PDone ;
    input [15:0]OuterAddress ;
    input [3:0]ResultIn ;
    input CLK ;
    input LP ;
    input INTR ;
    input CNNIMGLOAD ;
    input Rst ;
    inout EnableReadingFromCPU ;
    inout DecompressionDone ;
    inout DecompressionDone1 ;
    inout DecompressionDone2 ;
    inout readenable ;
    input [15:0]DataBus ;
    inout [15:0]Address ;
    inout [255:0]DecompressedData ;
    inout [255:0]DecompressedData1 ;
    inout [255:0]DecompressedData2 ;
    inout EnableReadingFromCPU1 ;
    inout EnableReadingFromCPU2 ;
    inout loadingimg ;
    inout loadingCNN ;
    output PClk ;
    output [255:0]DataFromRam ;
    inout [3:0]Result ;
    inout Done ;
    output ProcessEnable ;

    wire i8_reset2, nx2, loadenable, nx8, nx14, nx22, nx28, nx32, nx44, nx46, 
         nx52, nx54, nx62, nx66, nx70, nx74, nx82, i8_read2, zed, 
         i8_counterout1_1, i8_reset1, nx98, i8_counterout1_7, nx102, nx104, 
         nx110, i8_counterout1_5, i8_counterout1_4, i8_counterout1_3, 
         i8_counterout1_2, nx3092, i8_counterout1_0, nx128, nx136, nx152, nx3093, 
         nx182, nx3095, nx206, nx3097, nx230, nx3099, nx254, nx268, nx278, nx282, 
         nx298, i8_nx74, nx314, nx316, nx330, nx340, nx356, nx360, nx362, 
         i8_counterout2_5, nx370, nx374, nx376, i8_counterout2_4, nx3100, 
         i8_counterout2_3, nx3101, i8_counterout2_2, nx3102, i8_counterout2_1, 
         i8_counterout2_0, nx396, nx408, nx424, nx444, nx458, nx464, 
         i8_counterout2_7, i8_counterout2_6, nx480, nx494, nx514, nx520, nx528, 
         nx532, nx536, nx3104, nx540, nx546, nx558, nx560, nx572, i8_loadenableD, 
         nx588, nx602, nx610, nx618, nx622, i7_tmp, i7_counterout1_7, i7_start, 
         nx638, i7_reset2, i7_read2, i7_counterout2_7, nx648, nx650, nx654, 
         i7_counterout2_6, i7_counterout2_5, nx3107, i7_counterout2_4, nx3109, 
         i7_counterout2_3, nx3111, i7_counterout2_2, i7_counterout2_1, 
         i7_counterout2_0, nx674, nx690, nx708, nx724, nx740, nx758, nx772, 
         nx796, nx802, nx808, nx812, nx814, NOT_nx814, nx818, nx830, nx836, 
         i7_loadenableD, nx846, nx856, i7_counterout1_6, nx862, nx874, 
         i7_counterout1_5, nx3115, i7_counterout1_4, nx3116, nx894, 
         i7_counterout1_3, nx3117, nx912, i7_counterout1_2, nx3118, nx926, 
         i7_counterout1_1, nx940, i7_counterout1_0, nx952, nx960, nx974, nx994, 
         nx1014, nx1034, nx1054, nx1058, nx1078, nx1082, nx1084, nx1100, nx1110, 
         nx1128, nx1130, nx1134, nx1138, nx1140, nx1148, nx1154, nx1158, nx1174, 
         nx1176, nx1186, nx1188, nx1192, nx1202, nx1206, nx1216, nx1220, nx1230, 
         nx1234, nx1244, nx1248, nx1258, nx1262, nx1272, nx1276, nx1286, nx1290, 
         nx1300, nx1304, nx1314, nx1318, nx1328, nx1332, nx1342, nx1346, nx1356, 
         nx1360, nx1370, nx1374, nx1386, nx1388, nx1394, nx1398, nx1410, nx1422, 
         nx1434, nx1446, nx1458, nx1470, nx1482, nx1494, nx1506, nx1518, nx1530, 
         nx1542, nx1554, i5_MARo_0, i5_FAEN, nx1566, nx1576, nx1598, nx1604, 
         nx1606, nx1614, nx1616, nx1626, nx1634, nx1642, i5_MARo_1, nx1660, 
         nx1668, nx1670, i5_MARo_2, nx1682, nx1688, nx1696, nx1698, i5_MARo_3, 
         nx1708, nx1716, nx1724, nx1726, i5_MARo_4, nx1736, nx1744, nx1752, 
         nx1754, i5_MARo_5, nx1764, nx1772, nx1780, nx1782, i5_MARo_6, nx1794, 
         nx1800, nx1808, nx1810, i5_MARo_7, nx1820, nx1828, nx1836, nx1838, 
         i5_MARo_8, nx1848, nx1856, nx1864, nx1866, i5_MARo_9, nx1876, nx1884, 
         nx1892, nx1894, i5_MARo_10, nx1906, nx1912, nx1920, nx1922, i5_MARo_11, 
         nx1932, nx1940, nx1948, nx1950, i5_MARo_12, nx1960, nx1968, nx1976, 
         nx1978, i5_MARo_13, nx1988, nx1996, nx2004, nx2006, i5_MARo_14, nx2018, 
         nx2024, nx2032, nx2034, i5_MARo_15, nx2044, nx2052, nx2060, nx2062, 
         nx2068, nx2072, nx2080, nx2086, nx2098, nx2106, nx2108, nx2118, nx2122, 
         nx2134, nx2148, nx2160, nx2174, nx2186, nx2200, nx2212, nx2226, nx2238, 
         nx2252, nx2264, nx2278, nx2290, nx2304, nx2320, nx2334, nx2358, nx2382, 
         nx2406, nx2430, nx2444, nx2494, nx2512, nx2514, nx2520, nx2524, nx2548, 
         nx2572, nx2596, nx2620, nx2644, nx2668, nx2692, nx2708, nx2722, nx2746, 
         nx2770, nx2794, nx2818, nx2832, nx2880, nx2888, nx2902, nx2904, nx2910, 
         nx2914, nx2938, nx2962, nx2986, nx3010, nx3034, nx3058, nx3082, nx3098, 
         nx3112, nx3136, nx3160, nx3184, nx3208, nx3222, nx3272, nx3290, nx3292, 
         nx3298, nx3302, nx3326, nx3350, nx3374, nx3398, nx3422, nx3446, nx3470, 
         nx3486, nx3500, nx3524, nx3548, nx3572, nx3596, nx3610, nx3660, nx3668, 
         nx3682, nx3686, nx3688, nx3698, nx3702, nx3726, nx3750, nx3774, nx3798, 
         nx3822, nx3846, nx3870, nx3886, nx3900, nx3924, nx3948, nx3972, nx3996, 
         nx4010, nx4060, nx4074, nx4076, nx4082, nx4086, nx4110, nx4134, nx4158, 
         nx4182, nx4206, nx4230, nx4254, nx4270, nx4284, nx4308, nx4332, nx4356, 
         nx4380, nx4394, nx4446, nx4454, nx4468, nx4470, nx4476, nx4480, nx4504, 
         nx4528, nx4552, nx4576, nx4600, nx4624, nx4648, nx4664, nx4678, nx4702, 
         nx4726, nx4750, nx4774, nx4788, nx4838, nx4852, nx4854, nx4860, nx4864, 
         nx4888, nx4912, nx4936, nx4960, nx4984, nx5008, nx5032, nx5048, nx5062, 
         nx5086, nx5110, nx5134, nx5158, nx5172, nx5220, nx5228, nx5242, nx5246, 
         nx5248, nx5258, nx5262, nx5286, nx5310, nx5334, nx5358, nx5382, nx5406, 
         nx5430, nx5446, nx5460, nx5484, nx5508, nx5532, nx5556, nx5570, nx5620, 
         nx5634, nx5636, nx5642, nx5646, nx5670, nx5694, nx5718, nx5742, nx5766, 
         nx5790, nx5814, nx5830, nx5844, nx5868, nx5892, nx5916, nx5940, nx5954, 
         nx6002, nx6010, nx6024, nx6026, nx6032, nx6036, nx6060, nx6084, nx6108, 
         nx6132, nx6156, nx6180, nx6204, nx6220, nx6234, nx6258, nx6282, nx6306, 
         nx6330, nx6344, nx6394, nx6408, nx6410, nx6416, nx6420, nx6444, nx6468, 
         nx6492, nx6516, nx6540, nx6564, nx6588, nx6604, nx6618, nx6642, nx6666, 
         nx6690, nx6714, nx6728, nx6778, nx6786, nx6800, nx6802, nx6808, nx6812, 
         nx6836, nx6860, nx6884, nx6908, nx6932, nx6956, nx6980, nx6996, nx7010, 
         nx7034, nx7058, nx7082, nx7106, nx7120, nx7170, nx7184, nx7186, nx7192, 
         nx7196, nx7220, nx7244, nx7268, nx7292, nx7316, nx7340, nx7364, nx7380, 
         nx7394, nx7418, nx7442, nx7466, nx7490, nx7504, nx3127, nx3137, nx3147, 
         nx3157, nx3167, nx3177, nx3187, nx3197, nx3207, nx3217, nx3223, nx3225, 
         nx3227, nx3233, nx3235, nx3237, nx3247, nx3257, nx3267, nx3277, nx3283, 
         nx3293, nx3307, nx3317, nx3327, nx3337, nx3347, nx3357, nx3367, nx3377, 
         nx3383, nx3393, nx3407, nx3417, nx3427, nx3437, nx3447, nx3457, nx3467, 
         nx3477, nx3483, nx3493, nx3503, nx3518, nx3521, nx3523, nx3527, nx3533, 
         nx3537, nx3541, nx3545, nx3553, nx3555, nx3557, nx3561, nx3563, nx3565, 
         nx3569, nx3571, nx3575, nx3895, nx3899, nx3904, nx3907, nx3909, nx3917, 
         nx3919, nx3921, nx3925, nx3928, nx3930, nx3935, nx3938, nx3940, nx3943, 
         nx3947, nx3955, nx3959, nx3962, nx3967, nx3969, nx3971, nx3976, nx3979, 
         nx3985, nx3988, nx3993, nx3999, nx4002, nx4007, nx4011, nx4013, nx4016, 
         nx4019, nx4022, nx4026, nx4029, nx4033, nx4037, nx4041, nx4045, nx4050, 
         nx4053, nx4059, nx4063, nx4066, nx4073, nx4075, nx4079, nx4083, nx4090, 
         nx4093, nx4100, nx4107, nx4111, nx4114, nx4119, nx4124, nx4126, nx4131, 
         nx4138, nx4141, nx4148, nx4151, nx4155, nx4159, nx4162, nx4167, nx4171, 
         nx4177, nx4179, nx4181, nx4188, nx4191, nx4196, nx4198, nx4203, nx4207, 
         nx4209, nx4212, nx4215, nx4217, nx4220, nx4227, nx4231, nx4233, nx4237, 
         nx4239, nx4243, nx4246, nx4251, nx4255, nx4258, nx4261, nx4263, nx4267, 
         nx4271, nx4274, nx4277, nx4281, nx4283, nx4287, nx4293, nx4298, nx4301, 
         nx4303, nx4307, nx4309, nx4312, nx4315, nx4317, nx4318, nx4322, nx4327, 
         nx4331, nx4333, nx4336, nx4343, nx4345, nx4348, nx4353, nx4355, nx4359, 
         nx4367, nx4370, nx4374, nx4377, nx4379, nx4381, nx4383, nx4386, nx4389, 
         nx4393, nx4397, nx4399, nx4403, nx4405, nx4407, nx4409, nx4413, nx4417, 
         nx4419, nx4425, nx4427, nx4430, nx4434, nx4437, nx4441, nx4445, nx4447, 
         nx4453, nx4457, nx4460, nx4462, nx4465, nx4469, nx4475, nx4479, nx4485, 
         nx4487, nx4496, nx4501, nx4509, nx4511, nx4517, nx4522, nx4525, nx4532, 
         nx4535, nx4537, nx4542, nx4547, nx4553, nx4558, nx4565, nx4570, nx4577, 
         nx4582, nx4592, nx4613, nx4615, nx4618, nx4621, nx4625, nx4663, nx4665, 
         nx4668, nx4670, nx4673, nx4711, nx4715, nx4717, nx4720, nx4757, nx4759, 
         nx4763, nx4765, nx4804, nx4807, nx4809, nx4847, nx4851, nx4853, nx4894, 
         nx4897, nx4899, nx4937, nx4939, nx4942, nx4945, nx4985, nx4988, nx4990, 
         nx5029, nx5033, nx5035, nx5075, nx5078, nx5080, nx5119, nx5121, nx5124, 
         nx5126, nx5165, nx5169, nx5171, nx5209, nx5212, nx5215, nx5259, nx5263, 
         nx5266, nx5303, nx5305, nx5331, nx5333, nx5347, nx5349, nx5362, nx5375, 
         nx5389, nx5403, nx5415, nx5427, nx5441, nx5454, nx5467, nx5481, nx5497, 
         nx5509, nx5522, nx5535, nx5549, nx5562, nx5576, nx5589, nx5603, nx5615, 
         nx5628, nx5643, nx5659, nx5671, nx5684, nx5695, nx5697, nx5700, nx5703, 
         nx5707, nx5709, nx5712, nx5715, nx5719, nx5721, nx5724, nx5727, nx5731, 
         nx5733, nx5736, nx5739, nx5743, nx5745, nx5748, nx5751, nx5755, nx5757, 
         nx5760, nx5763, nx5767, nx5769, nx5772, nx5775, nx5779, nx5782, nx5785, 
         nx5787, nx5791, nx5793, nx5796, nx5799, nx5803, nx5805, nx5808, nx5811, 
         nx5815, nx5817, nx5820, nx5823, nx5827, nx5829, nx5833, nx5835, nx5838, 
         nx5841, nx5845, nx5847, nx5850, nx5853, nx5857, nx5859, nx5862, nx5865, 
         nx5869, nx5872, nx5875, nx5877, nx5881, nx5883, nx5886, nx5889, nx5893, 
         nx5895, nx5898, nx5901, nx5905, nx5907, nx5910, nx5913, nx5917, nx5919, 
         nx5922, nx5925, nx5929, nx5931, nx5934, nx5937, nx5941, nx5943, nx5946, 
         nx5949, nx5953, nx5955, nx5958, nx5961, nx5965, nx5967, nx5970, nx5973, 
         nx5977, nx5979, nx5982, nx5985, nx5989, nx5991, nx5994, nx5997, nx6001, 
         nx6003, nx6007, nx6009, nx6013, nx6015, nx6018, nx6021, nx6025, nx6027, 
         nx6031, nx6033, nx6037, nx6039, nx6042, nx6045, nx6049, nx6052, nx6055, 
         nx6057, nx6061, nx6063, nx6066, nx6069, nx6073, nx6075, nx6078, nx6081, 
         nx6085, nx6087, nx6090, nx6093, nx6097, nx6099, nx6102, nx6105, nx6109, 
         nx6111, nx6114, nx6117, nx6121, nx6123, nx6126, nx6129, nx6133, nx6135, 
         nx6138, nx6141, nx6145, nx6147, nx6150, nx6153, nx6157, nx6159, nx6162, 
         nx6165, nx6169, nx6171, nx6174, nx6177, nx6181, nx6183, nx6186, nx6189, 
         nx6193, nx6195, nx6198, nx6201, nx6205, nx6207, nx6210, nx6213, nx6217, 
         nx6219, nx6223, nx6225, nx6228, nx6231, nx6235, nx6237, nx6240, nx6243, 
         nx6247, nx6249, nx6252, nx6255, nx6259, nx6261, nx6264, nx6267, nx6271, 
         nx6273, nx6276, nx6279, nx6283, nx6285, nx6288, nx6291, nx6295, nx6297, 
         nx6300, nx6303, nx6307, nx6309, nx6312, nx6315, nx6319, nx6322, nx6325, 
         nx6327, nx6331, nx6333, nx6336, nx6339, nx6343, nx6345, nx6348, nx6350, 
         nx6353, nx6355, nx6358, nx6360, nx6363, nx6365, nx6368, nx6370, nx6373, 
         nx6375, nx6379, nx6381, nx6384, nx6387, nx6391, nx6393, nx6397, nx6399, 
         nx6402, nx6405, nx6409, nx6411, nx6415, nx6417, nx6421, nx6423, nx6426, 
         nx6429, nx6433, nx6435, nx6438, nx6441, nx6445, nx6447, nx6450, nx6453, 
         nx6457, nx6459, nx6462, nx6465, nx6469, nx6471, nx6474, nx6477, nx6481, 
         nx6483, nx6486, nx6489, nx6493, nx6496, nx6499, nx6501, nx6505, nx6507, 
         nx6510, nx6513, nx6517, nx6519, nx6522, nx6525, nx6529, nx6531, nx6534, 
         nx6537, nx6541, nx6543, nx6546, nx6549, nx6553, nx6555, nx6558, nx6561, 
         nx6565, nx6567, nx6570, nx6573, nx6577, nx6579, nx6582, nx6585, nx6589, 
         nx6591, nx6594, nx6597, nx6601, nx6603, nx6607, nx6609, nx6612, nx6615, 
         nx6619, nx6621, nx6624, nx6627, nx6631, nx6633, nx6636, nx6639, nx6643, 
         nx6645, nx6648, nx6651, nx6655, nx6657, nx6660, nx6663, nx6667, nx6669, 
         nx6672, nx6675, nx6679, nx6681, nx6684, nx6687, nx6691, nx6693, nx6696, 
         nx6699, nx6703, nx6705, nx6708, nx6711, nx6715, nx6717, nx6720, nx6723, 
         nx6727, nx6729, nx6732, nx6734, nx6737, nx6739, nx6742, nx6744, nx6747, 
         nx6749, nx6752, nx6754, nx6757, nx6761, nx6764, nx6766, nx6769, nx6771, 
         nx6775, nx6777, nx6781, nx6783, nx6787, nx6789, nx6792, nx6794, nx6797, 
         nx6799, nx6803, nx6805, nx6809, nx6811, nx6815, nx6817, nx6821, nx6823, 
         nx6826, nx6828, nx6831, nx6833, nx6837, nx6839, nx6842, nx6845, nx6849, 
         nx6851, nx6854, nx6857, nx6861, nx6863, nx6866, nx6869, nx6873, nx6875, 
         nx6878, nx6881, nx6885, nx6887, nx6890, nx6893, nx6897, nx6899, nx6902, 
         nx6905, nx6909, nx6911, nx6914, nx6917, nx6921, nx6923, nx6926, nx6929, 
         nx6933, nx6936, nx6939, nx6943, nx6946, nx6949, nx6953, nx6957, nx6960, 
         nx6963, nx6967, nx6970, nx6973, nx6977, nx6981, nx6984, nx6987, nx6991, 
         nx6995, nx6999, nx7002, nx7005, nx7009, nx7013, nx7016, nx7019, nx7023, 
         nx7026, nx7029, nx7033, nx7037, nx7039, nx7045, nx7048, nx7051, nx7057, 
         nx7063, nx7067, nx7072, nx7079, nx7081, nx7085, nx7088, nx7095, nx7098, 
         nx7100, nx7103, nx7107, nx7109, nx7115, nx7117, nx7121, nx7123, nx7126, 
         nx7129, nx7132, nx7137, nx7139, nx7143, nx7145, nx7148, nx7151, nx7157, 
         nx7159, nx7163, nx7165, nx7169, nx7173, nx7178, nx7181, nx7185, nx7189, 
         nx7197, nx7199, nx7202, nx7205, nx7209, nx7211, nx7214, nx7221, nx7223, 
         nx7226, nx7229, nx7233, nx7236, nx7241, nx7243, nx7247, nx7249, nx7253, 
         nx7257, nx7262, nx7265, nx7269, nx7272, nx7277, nx7279, nx7282, nx7284, 
         nx7287, nx7289, nx7293, nx7298, nx7301, nx7305, nx7307, nx7310, nx7313, 
         nx7319, nx7321, nx7325, nx7327, nx7330, nx7333, nx7339, nx7341, nx7344, 
         nx7347, nx7354, nx7356, nx7359, nx7361, nx7365, nx7367, nx7370, nx7377, 
         nx7381, nx7383, nx7390, nx7392, nx7395, nx7397, nx7399, nx7401, nx7403, 
         nx7405, nx7407, nx7409, nx7411, nx7413, nx7415, nx7417, nx7419, nx7421, 
         nx7423, nx7425, nx7427, nx7429, nx7431, nx7433, nx7435, nx7437, nx7439, 
         nx7441, nx7443, nx7445, nx7447, nx7449, nx7451, nx7455, nx7457, nx7459, 
         nx7461, nx7463, nx7465, nx7467, nx7469, nx7471, nx7473, nx7475, nx7477, 
         nx7479, nx7481, nx7483, nx7485, nx7487, nx7489, nx7491, nx7493, nx7495, 
         nx7497, nx7499, nx7501, nx7503, nx7505, nx7507, nx7509, nx7511, nx7515, 
         nx7517, nx7519, nx7521, nx7523, nx7525, nx7527, nx7529, nx7531, nx7537, 
         nx7539, nx7541, nx7551, nx7553, nx7555, nx7557, nx7559, nx7561, nx7563, 
         nx7565, nx7567, nx7569, nx7571, nx7575, nx7577, nx7579, nx7581, nx7583, 
         nx7587, nx7589, nx7591, nx7593, nx7595, nx7599, nx7601, nx7603, nx7605, 
         nx7607, nx7611, nx7613, nx7615, nx7617, nx7619, nx7623, nx7625, nx7627, 
         nx7629, nx7631, nx7633, nx7635, nx7637, nx7639, nx7643, nx7645, nx7647, 
         nx7649, nx7651, nx7655, nx7657, nx7659, nx7661, nx7663, nx7667, nx7669, 
         nx7671, nx7673, nx7675, nx7679, nx7681, nx7683, nx7685, nx7687, nx7691, 
         nx7693, nx7695, nx7697, nx7699, nx7703, nx7705, nx7707, nx7709, nx7711, 
         nx7715, nx7717, nx7719, nx7721, nx7723, nx7727, nx7729, nx7731, nx7733, 
         nx7735, nx7737, nx7739, nx7741, nx7743, nx7745, nx7747, nx7749, nx7751, 
         nx7753, nx7755, nx7757, nx7759, nx7761, nx7763, nx7765, nx7767, nx7769, 
         nx7771, nx7773, nx7775, nx7777, nx7779, nx7781, nx7783, nx7785, nx7787, 
         nx7789, nx7791, nx7793, nx7795, nx7797, nx7799, nx7801, nx7803, nx7805, 
         nx7807, nx7809, nx7811, nx7813, nx7815, nx7817, nx7819, nx7821, nx7823, 
         nx7825, nx7827, nx7829, nx7831, nx7833, nx7835, nx7837, nx7839, nx7841, 
         nx7843, nx7845, nx7847, nx7849, nx7851, nx7853, nx7855, nx7857, nx7859, 
         nx7861, nx7863, nx7865, nx7867, nx7869, nx7871, nx7873, nx7875, nx7877, 
         nx7879, nx7881, nx7883, nx7885, nx7887, nx7889, nx7891, nx7893, nx7895, 
         nx7897, nx7899, nx7901, nx7907, nx7909, nx7911, nx7913, nx7957, nx7959, 
         nx7961, nx8009, nx8011, nx8013, nx8015, nx8017, nx8019, nx8021, nx8023, 
         nx8025, nx8027, nx8029, nx8031, nx8033, nx8035, nx8037, nx8039, nx8041, 
         nx8043, nx8045, nx8047, nx8049, nx8051, nx8053, nx8055, nx8057, nx8059, 
         nx8061, nx8063, nx8065, nx8067, nx8069, nx8071, nx8073, nx8075, nx8077, 
         nx8079, nx8081, nx8083, nx8085, nx8087, nx8089, nx5, nx8093, nx8096, 
         nx8099, nx8102, nx8105, nx8108, nx8111, nx8114, nx8117, nx8120, nx8123, 
         nx8126, nx8129, nx8132, nx8135, nx8138, nx8141, nx8144, nx8147, nx8150, 
         nx8153, nx8156, nx8159, nx8162, nx8165, nx8168, nx8171, nx8174, nx8177, 
         nx8180, nx8183, nx8186, nx8189, nx8192, nx8195, nx8198, nx8201, nx8204, 
         nx8207, nx8210, nx8213, nx8216, nx8219, nx8222, nx8225, nx8228, nx8231, 
         nx8234, nx8237, nx8240, nx8243, nx8246, nx8249, nx8252, nx8255, nx8258, 
         nx8261, nx8264, nx8267, nx8270, nx8273, nx8276, nx8279, nx8282, nx8285, 
         nx8288, nx8291, nx8294, nx8297, nx8300, nx8303, nx8306, nx8309, nx8312, 
         nx8315, nx8318, nx8321, nx8324, nx8327, nx8330, nx8333, nx8336, nx8339, 
         nx8342, nx8345, nx8348, nx8351, nx8354, nx8357, nx8360, nx8363, nx8366, 
         nx8369, nx8372, nx8375, nx8378, nx8381, nx8384, nx8387, nx8390, nx8393, 
         nx8396, nx8399, nx8402, nx8405, nx8408, nx8411, nx8414, nx8417, nx8420, 
         nx8423, nx8426, nx8429, nx8432, nx8435, nx8438, nx8441, nx8444, nx8447, 
         nx8450, nx8453, nx8456, nx8459, nx8462, nx8465, nx8468, nx8471, nx8474, 
         nx8477, nx8480, nx8483, nx8486, nx8489, nx8492, nx8495, nx8498, nx8501, 
         nx8504, nx8507, nx8510, nx8513, nx8516, nx8519, nx8522, nx8525, nx8528, 
         nx8531, nx8534, nx8537, nx8540, nx8543, nx8546, nx8549, nx8552, nx8555, 
         nx8558, nx8561, nx8564, nx8567, nx8570, nx8573, nx8576, nx8579, nx8582, 
         nx8585, nx8588, nx8591, nx8594, nx8597, nx8600, nx8603, nx8606, nx8609, 
         nx8612, nx8615, nx8618, nx8621, nx8624, nx8627, nx8630, nx8633, nx8636, 
         nx8639, nx8642, nx8645, nx8648, nx8651, nx8654, nx8657, nx8660, nx8663, 
         nx8666, nx8669, nx8672, nx8675, nx8678, nx8681, nx8684, nx8687, nx8690, 
         nx8693, nx8696, nx8699, nx8702, nx8705, nx8708, nx8711, nx8714, nx8717, 
         nx8720, nx8723, nx8726, nx8729, nx8732, nx8735, nx8738, nx8741, nx8744, 
         nx8747, nx8750, nx8753, nx8756, nx8759, nx8762, nx8765, nx8768, nx8771, 
         nx8774, nx8777, nx8780, nx8783, nx8786, nx8789, nx8792, nx8795, nx8798, 
         nx8801, nx8804, nx8807, nx8810, nx8813, nx8816, nx8819, nx8822, nx8825, 
         nx8828, nx8831, nx8834, nx8837, nx8840, nx8843, nx8846, nx8849, nx8852, 
         nx8855, nx8858, nx8861, nx8864, nx8867, nx8870, nx8873, nx8876, nx8879, 
         nx8882, nx8885, nx8888, nx8891, nx8894, nx8897, nx8900, nx8903, nx8906, 
         nx8909, nx8912, nx8915, nx8918, nx8921, nx8924, nx8927, nx8930, nx8933, 
         nx8936, nx8939, nx8942, nx8945, nx8948, nx8951, nx8954, nx8957, nx8960, 
         nx8963, nx8966, nx8969, nx8972, nx8975, nx8978, nx8981, nx8984, nx8987, 
         nx8990, nx8993, nx8996, nx8999, nx9002, nx9005, nx9008, nx9011, nx9014, 
         nx9017, nx9020, nx9023, nx9026, nx9029, nx9032, nx9035, nx9038, nx9041, 
         nx9044, nx9047, nx9050, nx9053, nx9056, nx9059, nx9062, nx9065, nx9068, 
         nx9071, nx9074, nx9077, nx9080, nx9083, nx9086, nx9089, nx9092, nx9095, 
         nx9098, nx9101, nx9104, nx9107, nx9110, nx9113, nx9116, nx9119, nx9122, 
         nx9125, nx9128, nx9131, nx9134, nx9137, nx9140, nx9143, nx9146, nx9149, 
         nx9152, nx9155, nx9158, nx9161, nx9164, nx9167, nx9170, nx9173, nx9176, 
         nx9179, nx9182, nx9185, nx9188, nx9191, nx9194, nx9197, nx9200, nx9203, 
         nx9206, nx9209, nx9212, nx9215, nx9218, nx9221, nx9224, nx9227, nx9230, 
         nx9233, nx9236, nx9239, nx9242, nx9245, nx9248, nx9251, nx9254, nx9257, 
         nx9260, nx9263, nx9266, nx9269, nx9272, nx9274, nx9276, nx9278, nx9280, 
         nx9282, nx9284, nx9286, nx9288, nx9290, nx9292, nx9294, nx9296, nx9298, 
         nx9300, nx9302, nx9304, nx9306, nx9308, nx9310, nx9312, nx9314, nx9316, 
         nx9318, nx9320, nx9322, nx9324, nx9326, nx9328, nx9330, nx9332, nx9334, 
         nx9336, nx9338, nx9340, nx9342, nx9344, nx9346, nx9348, nx9350, nx9352, 
         nx9354, nx9356, nx9358, nx9360, nx9362, nx9364, nx9366, nx9368, nx9370, 
         nx9372, nx9374, nx9376, nx9378, nx9380, nx9382, nx9384, nx9386, nx9388, 
         nx9390, nx9392, nx9394, nx9396, nx9398, nx9400, nx9402, nx9404, nx9406, 
         nx9408;
    wire [10:0] \$dummy ;




    assign Result[3] = ResultIn[3] ;
    assign Result[2] = ResultIn[2] ;
    assign Result[1] = ResultIn[1] ;
    assign Result[0] = ResultIn[0] ;
    assign DecompressedData[254] = DecompressedData[255] ;
    assign DecompressedData[253] = DecompressedData[255] ;
    assign DecompressedData[238] = DecompressedData[239] ;
    assign DecompressedData[237] = DecompressedData[239] ;
    assign DecompressedData1[254] = DecompressedData1[255] ;
    assign DecompressedData1[253] = DecompressedData1[255] ;
    assign DecompressedData1[252] = DecompressedData1[255] ;
    assign DecompressedData1[251] = DecompressedData1[255] ;
    assign DecompressedData1[250] = DecompressedData1[255] ;
    assign DecompressedData1[249] = DecompressedData1[255] ;
    assign DecompressedData1[248] = DecompressedData1[255] ;
    assign DecompressedData1[247] = DecompressedData1[255] ;
    assign DecompressedData1[246] = DecompressedData1[255] ;
    assign DecompressedData1[245] = DecompressedData1[255] ;
    assign DecompressedData1[244] = DecompressedData1[255] ;
    assign DecompressedData1[243] = DecompressedData1[255] ;
    assign DecompressedData1[242] = DecompressedData1[255] ;
    assign DecompressedData1[241] = DecompressedData1[255] ;
    assign DecompressedData1[240] = DecompressedData1[255] ;
    assign DecompressedData1[239] = DecompressedData1[255] ;
    assign DecompressedData1[238] = DecompressedData1[255] ;
    assign DecompressedData1[237] = DecompressedData1[255] ;
    assign DecompressedData1[236] = DecompressedData1[255] ;
    assign DecompressedData1[235] = DecompressedData1[255] ;
    assign DecompressedData1[234] = DecompressedData1[255] ;
    assign DecompressedData1[233] = DecompressedData1[255] ;
    assign DecompressedData1[232] = DecompressedData1[255] ;
    assign DecompressedData1[231] = DecompressedData1[255] ;
    assign DecompressedData1[230] = DecompressedData1[255] ;
    assign DecompressedData1[229] = DecompressedData1[255] ;
    assign DecompressedData1[228] = DecompressedData1[255] ;
    assign DecompressedData1[227] = DecompressedData1[255] ;
    assign DecompressedData1[226] = DecompressedData1[255] ;
    assign DecompressedData1[225] = DecompressedData1[255] ;
    assign DecompressedData1[224] = DecompressedData1[255] ;
    assign DecompressedData2[254] = DecompressedData2[255] ;
    assign DecompressedData2[253] = DecompressedData2[255] ;
    assign DecompressedData2[238] = DecompressedData2[239] ;
    assign DecompressedData2[237] = DecompressedData2[239] ;
    assign DecompressedData2[222] = DecompressedData2[223] ;
    assign DecompressedData2[221] = DecompressedData2[223] ;
    assign DecompressedData2[206] = DecompressedData2[207] ;
    assign DecompressedData2[205] = DecompressedData2[207] ;
    assign DecompressedData2[190] = DecompressedData2[191] ;
    assign DecompressedData2[189] = DecompressedData2[191] ;
    assign DecompressedData2[174] = DecompressedData2[175] ;
    assign DecompressedData2[173] = DecompressedData2[175] ;
    assign DecompressedData2[158] = DecompressedData2[159] ;
    assign DecompressedData2[157] = DecompressedData2[159] ;
    assign DecompressedData2[142] = DecompressedData2[143] ;
    assign DecompressedData2[141] = DecompressedData2[143] ;
    assign DecompressedData2[126] = DecompressedData2[127] ;
    assign DecompressedData2[125] = DecompressedData2[127] ;
    assign DecompressedData2[110] = DecompressedData2[111] ;
    assign DecompressedData2[109] = DecompressedData2[111] ;
    assign DecompressedData2[94] = DecompressedData2[95] ;
    assign DecompressedData2[93] = DecompressedData2[95] ;
    assign DecompressedData2[78] = DecompressedData2[79] ;
    assign DecompressedData2[77] = DecompressedData2[79] ;
    assign DecompressedData2[62] = DecompressedData2[63] ;
    assign DecompressedData2[61] = DecompressedData2[63] ;
    assign DecompressedData2[46] = DecompressedData2[47] ;
    assign DecompressedData2[45] = DecompressedData2[47] ;
    assign DecompressedData2[30] = DecompressedData2[31] ;
    assign DecompressedData2[29] = DecompressedData2[31] ;
    assign DecompressedData2[14] = DecompressedData2[15] ;
    assign DecompressedData2[13] = DecompressedData2[15] ;
    assign PClk = CLK ;
    fake_vcc ix3 (.Y (nx2)) ;
    fake_gnd ix2589 (.Y (DecompressedData1[255])) ;
    nor02_2x ix631 (.Y (loadingimg), .A0 (CNNIMGLOAD), .A1 (nx7957)) ;
    nor02_2x ix83 (.Y (nx82), .A0 (LP), .A1 (nx3518)) ;
    nor02_2x ix3519 (.Y (nx3518), .A0 (nx74), .A1 (nx7737)) ;
    nor02_2x ix75 (.Y (nx74), .A0 (nx3521), .A1 (Rst)) ;
    inv01 ix3522 (.Y (nx3521), .A (INTR)) ;
    nor02_2x ix67 (.Y (nx66), .A0 (nx3527), .A1 (nx3533)) ;
    nand04 ix3528 (.Y (nx3527), .A0 (nx8), .A1 (nx14), .A2 (nx22), .A3 (nx28)) ;
    nor02_2x ix9 (.Y (nx8), .A0 (DataBus[8]), .A1 (DataBus[9])) ;
    nor02_2x ix15 (.Y (nx14), .A0 (DataBus[10]), .A1 (DataBus[11])) ;
    nor02_2x ix23 (.Y (nx22), .A0 (DataBus[12]), .A1 (DataBus[13])) ;
    nor02_2x ix29 (.Y (nx28), .A0 (DataBus[0]), .A1 (DataBus[1])) ;
    nand04 ix3534 (.Y (nx3533), .A0 (nx46), .A1 (nx52), .A2 (nx3541), .A3 (
           nx7907)) ;
    nor03_2x ix47 (.Y (nx46), .A0 (DataBus[2]), .A1 (DataBus[3]), .A2 (nx3537)
             ) ;
    inv01 ix3538 (.Y (nx3537), .A (nx44)) ;
    nor02_2x ix45 (.Y (nx44), .A0 (DataBus[4]), .A1 (DataBus[5])) ;
    nor02_2x ix53 (.Y (nx52), .A0 (DataBus[6]), .A1 (DataBus[7])) ;
    nor02_2x ix3542 (.Y (nx3541), .A0 (DataBus[14]), .A1 (DataBus[15])) ;
    dff i1_L_reg_Q (.Q (loadenable), .QB (\$dummy [0]), .D (nx82), .CLK (nx70)
        ) ;
    nand02 ix71 (.Y (nx70), .A0 (nx7737), .A1 (nx3521)) ;
    inv01 ix3546 (.Y (nx3545), .A (Rst)) ;
    nor02_2x ix91 (.Y (loadingCNN), .A0 (nx7741), .A1 (nx7957)) ;
    dff i0_L_reg_Q (.Q (ProcessEnable), .QB (nx3563), .D (nx1576), .CLK (nx1566)
        ) ;
    nor02_2x ix1577 (.Y (nx1576), .A0 (nx3553), .A1 (nx3557)) ;
    nor02_2x ix3554 (.Y (nx3553), .A0 (nx3555), .A1 (INTR)) ;
    inv01 ix3556 (.Y (nx3555), .A (PDone)) ;
    nand02 ix3558 (.Y (nx3557), .A0 (LP), .A1 (nx3545)) ;
    nand02 ix1567 (.Y (nx1566), .A0 (nx3561), .A1 (nx3545)) ;
    nor02_2x ix3562 (.Y (nx3561), .A0 (PDone), .A1 (INTR)) ;
    nand02 ix7553 (.Y (Done), .A0 (nx3565), .A1 (nx3555)) ;
    nand03 ix3566 (.Y (nx3565), .A0 (nx32), .A1 (nx46), .A2 (nx62)) ;
    nor02_2x ix33 (.Y (nx32), .A0 (nx3569), .A1 (nx3571)) ;
    nand02 ix3570 (.Y (nx3569), .A0 (nx8), .A1 (nx14)) ;
    nand02 ix3572 (.Y (nx3571), .A0 (nx22), .A1 (nx28)) ;
    nor03_2x ix63 (.Y (nx62), .A0 (DataBus[6]), .A1 (DataBus[7]), .A2 (nx3575)
             ) ;
    nand02 ix3576 (.Y (nx3575), .A0 (nx3541), .A1 (nx7907)) ;
    tri01 tri_DataFromRam_0 (.Y (DataFromRam[0]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_1 (.Y (DataFromRam[1]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_2 (.Y (DataFromRam[2]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_3 (.Y (DataFromRam[3]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_4 (.Y (DataFromRam[4]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_5 (.Y (DataFromRam[5]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_6 (.Y (DataFromRam[6]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_7 (.Y (DataFromRam[7]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_8 (.Y (DataFromRam[8]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_9 (.Y (DataFromRam[9]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_10 (.Y (DataFromRam[10]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_11 (.Y (DataFromRam[11]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_12 (.Y (DataFromRam[12]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_13 (.Y (DataFromRam[13]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_14 (.Y (DataFromRam[14]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_15 (.Y (DataFromRam[15]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_16 (.Y (DataFromRam[16]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_17 (.Y (DataFromRam[17]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_18 (.Y (DataFromRam[18]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_19 (.Y (DataFromRam[19]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_20 (.Y (DataFromRam[20]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_21 (.Y (DataFromRam[21]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_22 (.Y (DataFromRam[22]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_23 (.Y (DataFromRam[23]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_24 (.Y (DataFromRam[24]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_25 (.Y (DataFromRam[25]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_26 (.Y (DataFromRam[26]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_27 (.Y (DataFromRam[27]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_28 (.Y (DataFromRam[28]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_29 (.Y (DataFromRam[29]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_30 (.Y (DataFromRam[30]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_31 (.Y (DataFromRam[31]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_32 (.Y (DataFromRam[32]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_33 (.Y (DataFromRam[33]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_34 (.Y (DataFromRam[34]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_35 (.Y (DataFromRam[35]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_36 (.Y (DataFromRam[36]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_37 (.Y (DataFromRam[37]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_38 (.Y (DataFromRam[38]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_39 (.Y (DataFromRam[39]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_40 (.Y (DataFromRam[40]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_41 (.Y (DataFromRam[41]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_42 (.Y (DataFromRam[42]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_43 (.Y (DataFromRam[43]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_44 (.Y (DataFromRam[44]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_45 (.Y (DataFromRam[45]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_46 (.Y (DataFromRam[46]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_47 (.Y (DataFromRam[47]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_48 (.Y (DataFromRam[48]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_49 (.Y (DataFromRam[49]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_50 (.Y (DataFromRam[50]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_51 (.Y (DataFromRam[51]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_52 (.Y (DataFromRam[52]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_53 (.Y (DataFromRam[53]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_54 (.Y (DataFromRam[54]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_55 (.Y (DataFromRam[55]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_56 (.Y (DataFromRam[56]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_57 (.Y (DataFromRam[57]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_58 (.Y (DataFromRam[58]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_59 (.Y (DataFromRam[59]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_60 (.Y (DataFromRam[60]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_61 (.Y (DataFromRam[61]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_62 (.Y (DataFromRam[62]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_63 (.Y (DataFromRam[63]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_64 (.Y (DataFromRam[64]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_65 (.Y (DataFromRam[65]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_66 (.Y (DataFromRam[66]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_67 (.Y (DataFromRam[67]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_68 (.Y (DataFromRam[68]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_69 (.Y (DataFromRam[69]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_70 (.Y (DataFromRam[70]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_71 (.Y (DataFromRam[71]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_72 (.Y (DataFromRam[72]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_73 (.Y (DataFromRam[73]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_74 (.Y (DataFromRam[74]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_75 (.Y (DataFromRam[75]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_76 (.Y (DataFromRam[76]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_77 (.Y (DataFromRam[77]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_78 (.Y (DataFromRam[78]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_79 (.Y (DataFromRam[79]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_80 (.Y (DataFromRam[80]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_81 (.Y (DataFromRam[81]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_82 (.Y (DataFromRam[82]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_83 (.Y (DataFromRam[83]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_84 (.Y (DataFromRam[84]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_85 (.Y (DataFromRam[85]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_86 (.Y (DataFromRam[86]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_87 (.Y (DataFromRam[87]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_88 (.Y (DataFromRam[88]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_89 (.Y (DataFromRam[89]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_90 (.Y (DataFromRam[90]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_91 (.Y (DataFromRam[91]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_92 (.Y (DataFromRam[92]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_93 (.Y (DataFromRam[93]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_94 (.Y (DataFromRam[94]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_95 (.Y (DataFromRam[95]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_96 (.Y (DataFromRam[96]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_97 (.Y (DataFromRam[97]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_98 (.Y (DataFromRam[98]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_99 (.Y (DataFromRam[99]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_100 (.Y (DataFromRam[100]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_101 (.Y (DataFromRam[101]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_102 (.Y (DataFromRam[102]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_103 (.Y (DataFromRam[103]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_104 (.Y (DataFromRam[104]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_105 (.Y (DataFromRam[105]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_106 (.Y (DataFromRam[106]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_107 (.Y (DataFromRam[107]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_108 (.Y (DataFromRam[108]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_109 (.Y (DataFromRam[109]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_110 (.Y (DataFromRam[110]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_111 (.Y (DataFromRam[111]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_112 (.Y (DataFromRam[112]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_113 (.Y (DataFromRam[113]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_114 (.Y (DataFromRam[114]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_115 (.Y (DataFromRam[115]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_116 (.Y (DataFromRam[116]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_117 (.Y (DataFromRam[117]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_118 (.Y (DataFromRam[118]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_119 (.Y (DataFromRam[119]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_120 (.Y (DataFromRam[120]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_121 (.Y (DataFromRam[121]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_122 (.Y (DataFromRam[122]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_123 (.Y (DataFromRam[123]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_124 (.Y (DataFromRam[124]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_125 (.Y (DataFromRam[125]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_126 (.Y (DataFromRam[126]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_127 (.Y (DataFromRam[127]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_128 (.Y (DataFromRam[128]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_129 (.Y (DataFromRam[129]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_130 (.Y (DataFromRam[130]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_131 (.Y (DataFromRam[131]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_132 (.Y (DataFromRam[132]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_133 (.Y (DataFromRam[133]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_134 (.Y (DataFromRam[134]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_135 (.Y (DataFromRam[135]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_136 (.Y (DataFromRam[136]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_137 (.Y (DataFromRam[137]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_138 (.Y (DataFromRam[138]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_139 (.Y (DataFromRam[139]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_140 (.Y (DataFromRam[140]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_141 (.Y (DataFromRam[141]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_142 (.Y (DataFromRam[142]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_143 (.Y (DataFromRam[143]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_144 (.Y (DataFromRam[144]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_145 (.Y (DataFromRam[145]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_146 (.Y (DataFromRam[146]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_147 (.Y (DataFromRam[147]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_148 (.Y (DataFromRam[148]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_149 (.Y (DataFromRam[149]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_150 (.Y (DataFromRam[150]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_151 (.Y (DataFromRam[151]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_152 (.Y (DataFromRam[152]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_153 (.Y (DataFromRam[153]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_154 (.Y (DataFromRam[154]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_155 (.Y (DataFromRam[155]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_156 (.Y (DataFromRam[156]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_157 (.Y (DataFromRam[157]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_158 (.Y (DataFromRam[158]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_159 (.Y (DataFromRam[159]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_160 (.Y (DataFromRam[160]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_161 (.Y (DataFromRam[161]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_162 (.Y (DataFromRam[162]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_163 (.Y (DataFromRam[163]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_164 (.Y (DataFromRam[164]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_165 (.Y (DataFromRam[165]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_166 (.Y (DataFromRam[166]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_167 (.Y (DataFromRam[167]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_168 (.Y (DataFromRam[168]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_169 (.Y (DataFromRam[169]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_170 (.Y (DataFromRam[170]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_171 (.Y (DataFromRam[171]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_172 (.Y (DataFromRam[172]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_173 (.Y (DataFromRam[173]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_174 (.Y (DataFromRam[174]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_175 (.Y (DataFromRam[175]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_176 (.Y (DataFromRam[176]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_177 (.Y (DataFromRam[177]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_178 (.Y (DataFromRam[178]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_179 (.Y (DataFromRam[179]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_180 (.Y (DataFromRam[180]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_181 (.Y (DataFromRam[181]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_182 (.Y (DataFromRam[182]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_183 (.Y (DataFromRam[183]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_184 (.Y (DataFromRam[184]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_185 (.Y (DataFromRam[185]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_186 (.Y (DataFromRam[186]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_187 (.Y (DataFromRam[187]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_188 (.Y (DataFromRam[188]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_189 (.Y (DataFromRam[189]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_190 (.Y (DataFromRam[190]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_191 (.Y (DataFromRam[191]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_192 (.Y (DataFromRam[192]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_193 (.Y (DataFromRam[193]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_194 (.Y (DataFromRam[194]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_195 (.Y (DataFromRam[195]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_196 (.Y (DataFromRam[196]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_197 (.Y (DataFromRam[197]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_198 (.Y (DataFromRam[198]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_199 (.Y (DataFromRam[199]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_200 (.Y (DataFromRam[200]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_201 (.Y (DataFromRam[201]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_202 (.Y (DataFromRam[202]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_203 (.Y (DataFromRam[203]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_204 (.Y (DataFromRam[204]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_205 (.Y (DataFromRam[205]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_206 (.Y (DataFromRam[206]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_207 (.Y (DataFromRam[207]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_208 (.Y (DataFromRam[208]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_209 (.Y (DataFromRam[209]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_210 (.Y (DataFromRam[210]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_211 (.Y (DataFromRam[211]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_212 (.Y (DataFromRam[212]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_213 (.Y (DataFromRam[213]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_214 (.Y (DataFromRam[214]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_215 (.Y (DataFromRam[215]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_216 (.Y (DataFromRam[216]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_217 (.Y (DataFromRam[217]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_218 (.Y (DataFromRam[218]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_219 (.Y (DataFromRam[219]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_220 (.Y (DataFromRam[220]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_221 (.Y (DataFromRam[221]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_222 (.Y (DataFromRam[222]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_223 (.Y (DataFromRam[223]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_224 (.Y (DataFromRam[224]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_225 (.Y (DataFromRam[225]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_226 (.Y (DataFromRam[226]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_227 (.Y (DataFromRam[227]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_228 (.Y (DataFromRam[228]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_229 (.Y (DataFromRam[229]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_230 (.Y (DataFromRam[230]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_231 (.Y (DataFromRam[231]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_232 (.Y (DataFromRam[232]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_233 (.Y (DataFromRam[233]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_234 (.Y (DataFromRam[234]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_235 (.Y (DataFromRam[235]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_236 (.Y (DataFromRam[236]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_237 (.Y (DataFromRam[237]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_238 (.Y (DataFromRam[238]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_239 (.Y (DataFromRam[239]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_240 (.Y (DataFromRam[240]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_241 (.Y (DataFromRam[241]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_242 (.Y (DataFromRam[242]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_243 (.Y (DataFromRam[243]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_244 (.Y (DataFromRam[244]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_245 (.Y (DataFromRam[245]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_246 (.Y (DataFromRam[246]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_247 (.Y (DataFromRam[247]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_248 (.Y (DataFromRam[248]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_249 (.Y (DataFromRam[249]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_250 (.Y (DataFromRam[250]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_251 (.Y (DataFromRam[251]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_252 (.Y (DataFromRam[252]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_253 (.Y (DataFromRam[253]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_254 (.Y (DataFromRam[254]), .A (nx2), .E (
          DecompressedData1[255])) ;
    tri01 tri_DataFromRam_255 (.Y (DataFromRam[255]), .A (nx2), .E (
          DecompressedData1[255])) ;
    aoi21 ix611 (.Y (nx610), .A0 (nx7765), .A1 (zed), .B0 (nx4198)) ;
    nor02_2x ix3896 (.Y (nx3895), .A0 (nx3093), .A1 (nx282)) ;
    nand03 ix191 (.Y (nx3093), .A0 (nx3899), .A1 (nx4019), .A2 (nx4033)) ;
    nor02_2x ix3900 (.Y (nx3899), .A0 (i8_counterout1_0), .A1 (i8_counterout1_1)
             ) ;
    oai21 ix3128 (.Y (nx3127), .A0 (nx3904), .A1 (nx7805), .B0 (nx4196)) ;
    nor02_2x ix3905 (.Y (nx3904), .A0 (nx136), .A1 (nx128)) ;
    oai21 ix137 (.Y (nx136), .A0 (nx3907), .A1 (nx3909), .B0 (nx4188)) ;
    dff reg_i8_counterout1_0 (.Q (i8_counterout1_0), .QB (nx3907), .D (nx3127), 
        .CLK (CLK)) ;
    oai21 ix3910 (.Y (nx3909), .A0 (nx7741), .A1 (nx7401), .B0 (nx7769)) ;
    dffr i8_ix75 (.Q (i8_nx74), .QB (\$dummy [1]), .D (nx2), .CLK (CLK), .R (
         nx98)) ;
    nor02_2x ix99 (.Y (nx98), .A0 (nx3917), .A1 (nx3919)) ;
    nand02 ix3918 (.Y (nx3917), .A0 (CNNIMGLOAD), .A1 (nx7907)) ;
    nand02 ix3920 (.Y (nx3919), .A0 (nx7779), .A1 (nx4083)) ;
    dffs_ni i8_reg_start (.Q (\$dummy [2]), .QB (nx3921), .D (nx3293), .CLK (CLK
            ), .S (nx588)) ;
    nor02_2x ix3294 (.Y (nx3293), .A0 (nx7775), .A1 (nx3104)) ;
    nor02_2x ix579 (.Y (nx3104), .A0 (nx3925), .A1 (nx7769)) ;
    nor02_2x ix573 (.Y (nx572), .A0 (nx3917), .A1 (nx3928)) ;
    nand02 ix3929 (.Y (nx3928), .A0 (nx7775), .A1 (nx3930)) ;
    nor02_2x ix3284 (.Y (nx3283), .A0 (nx3930), .A1 (nx546)) ;
    nand03 ix547 (.Y (nx546), .A0 (nx3935), .A1 (nx4181), .A2 (nx3955)) ;
    nand03 ix529 (.Y (nx528), .A0 (nx7781), .A1 (nx7911), .A2 (i8_counterout2_3)
           ) ;
    nor02_2x ix3939 (.Y (nx3938), .A0 (nx3940), .A1 (nx4126)) ;
    oai21 ix3208 (.Y (nx3207), .A0 (nx3943), .A1 (nx7785), .B0 (nx4179)) ;
    nand02 ix377 (.Y (nx376), .A0 (nx3947), .A1 (nx7737)) ;
    nor02_2x ix3948 (.Y (nx3947), .A0 (i8_reset2), .A1 (nx7741)) ;
    dffr i8_ix97 (.Q (i8_reset2), .QB (nx3925), .D (nx2), .CLK (CLK), .R (nx572)
         ) ;
    dff reg_i8_counterout2_0 (.Q (i8_counterout2_0), .QB (nx3940), .D (nx3207), 
        .CLK (CLK)) ;
    nor02_2x ix537 (.Y (nx536), .A0 (nx3959), .A1 (nx4093)) ;
    nor02_2x ix3960 (.Y (nx3959), .A0 (nx360), .A1 (nx356)) ;
    nand04 ix361 (.Y (nx360), .A0 (nx3962), .A1 (nx3979), .A2 (nx4059), .A3 (
           i8_counterout1_0)) ;
    nor02_2x ix3963 (.Y (nx3962), .A0 (i8_counterout1_4), .A1 (i8_counterout1_5)
             ) ;
    oai22 ix207 (.Y (nx206), .A0 (nx3967), .A1 (nx3969), .B0 (nx3095), .B1 (
          nx104)) ;
    dff reg_i8_counterout1_4 (.Q (i8_counterout1_4), .QB (nx3967), .D (nx3157), 
        .CLK (CLK)) ;
    mux21 ix3970 (.Y (nx3969), .A0 (nx7769), .A1 (nx3093), .S0 (nx7801)) ;
    nor03_2x ix3972 (.Y (nx3971), .A0 (nx7415), .A1 (nx7741), .A2 (nx7401)) ;
    nand04 ix299 (.Y (nx298), .A0 (nx3976), .A1 (nx4083), .A2 (loadingCNN), .A3 (
           nx7775)) ;
    oai21 ix3977 (.Y (nx3976), .A0 (nx3093), .A1 (nx282), .B0 (nx3955)) ;
    nand03 ix283 (.Y (nx282), .A0 (nx3962), .A1 (nx3979), .A2 (nx4059)) ;
    oai22 ix255 (.Y (nx254), .A0 (nx3979), .A1 (nx3985), .B0 (nx3099), .B1 (
          nx104)) ;
    mux21 ix3986 (.Y (nx3985), .A0 (nx7769), .A1 (nx3097), .S0 (nx7801)) ;
    nand04 ix239 (.Y (nx3097), .A0 (nx3988), .A1 (nx4033), .A2 (nx3967), .A3 (
           nx4050)) ;
    nor03_2x ix3989 (.Y (nx3988), .A0 (i8_counterout1_0), .A1 (i8_counterout1_1)
             , .A2 (i8_counterout1_2)) ;
    oai21 ix3198 (.Y (nx3197), .A0 (nx3993), .A1 (nx7803), .B0 (nx4075)) ;
    aoi322 ix3994 (.Y (nx3993), .A0 (nx330), .A1 (nx54), .A2 (nx7413), .B0 (
           nx3899), .B1 (nx7799), .C0 (i8_counterout1_1), .C1 (nx340)) ;
    nand02 ix331 (.Y (nx330), .A0 (DataBus[14]), .A1 (DataBus[15])) ;
    inv01 ix55 (.Y (nx54), .A (nx3541)) ;
    mux21 ix341 (.Y (nx340), .A0 (nx7413), .A1 (nx3907), .S0 (nx7799)) ;
    nand02 ix4000 (.Y (nx3999), .A0 (loadingCNN), .A1 (nx316)) ;
    nand03 ix317 (.Y (nx316), .A0 (nx4002), .A1 (i8_read2), .A2 (nx7775)) ;
    nand02 ix4003 (.Y (nx4002), .A0 (nx7413), .A1 (zed)) ;
    nor03_2x ix541 (.Y (nx540), .A0 (nx4007), .A1 (nx3093), .A2 (nx282)) ;
    nand02 ix4008 (.Y (nx4007), .A0 (i8_reset2), .A1 (nx7413)) ;
    dffs_ni i8_reg_read2 (.Q (i8_read2), .QB (nx3930), .D (nx3283), .CLK (CLK), 
            .S (nx560)) ;
    nand03 ix561 (.Y (nx560), .A0 (nx546), .A1 (nx4011), .A2 (nx7775)) ;
    nand04 ix4012 (.Y (nx4011), .A0 (nx4013), .A1 (nx4045), .A2 (nx3541), .A3 (
           nx7395)) ;
    nand03 ix167 (.Y (nx3092), .A0 (nx3907), .A1 (nx4016), .A2 (nx4019)) ;
    dff reg_i8_counterout1_1 (.Q (i8_counterout1_1), .QB (nx4016), .D (nx3197), 
        .CLK (CLK)) ;
    oai21 ix3138 (.Y (nx3137), .A0 (nx4022), .A1 (nx7803), .B0 (nx4026)) ;
    aoi322 ix4023 (.Y (nx4022), .A0 (nx7413), .A1 (DataBus[15]), .A2 (
           DataBus[14]), .B0 (nx3988), .B1 (nx7799), .C0 (i8_counterout1_2), .C1 (
           nx152)) ;
    dff reg_i8_counterout1_2 (.Q (i8_counterout1_2), .QB (nx4019), .D (nx3137), 
        .CLK (CLK)) ;
    mux21 ix153 (.Y (nx152), .A0 (nx7413), .A1 (nx3899), .S0 (nx7799)) ;
    oai21 ix4027 (.Y (nx4026), .A0 (nx3917), .A1 (nx4029), .B0 (i8_counterout1_2
          )) ;
    oai21 ix315 (.Y (nx314), .A0 (nx7769), .A1 (nx3955), .B0 (i8_read2)) ;
    oai22 ix183 (.Y (nx182), .A0 (nx4033), .A1 (nx4037), .B0 (nx3093), .B1 (
          nx104)) ;
    mux21 ix4038 (.Y (nx4037), .A0 (nx7769), .A1 (nx3092), .S0 (nx7799)) ;
    nand02 ix105 (.Y (nx104), .A0 (nx4041), .A1 (nx7737)) ;
    nor02_2x ix4042 (.Y (nx4041), .A0 (nx7413), .A1 (nx7741)) ;
    dff reg_i8_counterout1_3 (.Q (i8_counterout1_3), .QB (nx4033), .D (nx3147), 
        .CLK (CLK)) ;
    nor03_2x ix4046 (.Y (nx4045), .A0 (i8_counterout1_4), .A1 (i8_counterout1_5)
             , .A2 (nx278)) ;
    oai22 ix231 (.Y (nx230), .A0 (nx4050), .A1 (nx4053), .B0 (nx3097), .B1 (
          nx104)) ;
    dff reg_i8_counterout1_5 (.Q (i8_counterout1_5), .QB (nx4050), .D (nx3167), 
        .CLK (CLK)) ;
    mux21 ix4054 (.Y (nx4053), .A0 (nx7769), .A1 (nx3095), .S0 (nx7799)) ;
    nand04 ix215 (.Y (nx3095), .A0 (nx3899), .A1 (nx4019), .A2 (nx4033), .A3 (
           nx3967)) ;
    nand02 ix279 (.Y (nx278), .A0 (nx3979), .A1 (nx4059)) ;
    oai21 ix3188 (.Y (nx3187), .A0 (nx4063), .A1 (nx7803), .B0 (nx4073)) ;
    nor02_2x ix4064 (.Y (nx4063), .A0 (nx268), .A1 (nx110)) ;
    nor02_2x ix269 (.Y (nx268), .A0 (nx4066), .A1 (nx104)) ;
    dff reg_i8_counterout1_7 (.Q (i8_counterout1_7), .QB (nx4059), .D (nx3187), 
        .CLK (CLK)) ;
    nor03_2x ix111 (.Y (nx110), .A0 (nx4059), .A1 (nx7415), .A2 (nx7799)) ;
    oai21 ix4074 (.Y (nx4073), .A0 (nx3917), .A1 (nx4029), .B0 (i8_counterout1_7
          )) ;
    oai21 ix4076 (.Y (nx4075), .A0 (nx3917), .A1 (nx4029), .B0 (i8_counterout1_1
          )) ;
    nand02 ix263 (.Y (nx3099), .A0 (nx4079), .A1 (nx3979)) ;
    dff i8_counterout1_6 (.Q (\$dummy [3]), .QB (nx3979), .D (nx3177), .CLK (CLK
        )) ;
    dffsr_ni i8_ix263 (.Q (EnableReadingFromCPU2), .QB (nx4083), .D (
             DecompressedData1[255]), .CLK (CLK), .S (nx610), .R (nx622)) ;
    nor02ii ix623 (.Y (nx622), .A0 (nx610), .A1 (nx618)) ;
    oai221 ix619 (.Y (nx618), .A0 (zed), .A1 (nx362), .B0 (DataBus[14]), .B1 (
           DataBus[15]), .C0 (nx7775)) ;
    nand04 ix363 (.Y (nx362), .A0 (nx4045), .A1 (i8_counterout1_0), .A2 (nx4090)
           , .A3 (nx4016)) ;
    nor02_2x ix4091 (.Y (nx4090), .A0 (i8_counterout1_2), .A1 (i8_counterout1_3)
             ) ;
    nand03 ix357 (.Y (nx356), .A0 (nx4019), .A1 (nx4033), .A2 (nx4016)) ;
    nor02_2x ix4094 (.Y (nx4093), .A0 (nx532), .A1 (nx514)) ;
    nand04 ix533 (.Y (nx532), .A0 (nx7781), .A1 (nx7911), .A2 (i8_counterout2_3)
           , .A3 (i8_counterout2_4)) ;
    inv01 ix3228 (.Y (nx3227), .A (nx4100)) ;
    nor02_2x ix4101 (.Y (nx4100), .A0 (nx3223), .A1 (nx3225)) ;
    nor02_2x ix3224 (.Y (nx3223), .A0 (nx7961), .A1 (nx7419)) ;
    dff reg_i8_counterout2_2 (.Q (i8_counterout2_2), .QB (\$dummy [4]), .D (
        nx3227), .CLK (CLK)) ;
    nand03 ix371 (.Y (nx370), .A0 (nx7811), .A1 (nx7395), .A2 (nx7777)) ;
    nand02 ix4108 (.Y (nx4107), .A0 (i8_reset2), .A1 (zed)) ;
    aoi32 ix3226 (.Y (nx3225), .A0 (nx7811), .A1 (nx7395), .A2 (nx7777), .B0 (
          nx4111), .B1 (nx3102)) ;
    nor03_2x ix4112 (.Y (nx4111), .A0 (nx408), .A1 (nx7427), .A2 (nx7401)) ;
    nor02_2x ix409 (.Y (nx408), .A0 (nx7961), .A1 (nx7813)) ;
    nor02_2x ix4115 (.Y (nx4114), .A0 (i8_counterout2_0), .A1 (i8_counterout2_1)
             ) ;
    dff reg_i8_counterout2_1 (.Q (i8_counterout2_1), .QB (nx4126), .D (nx3217), 
        .CLK (CLK)) ;
    oai21 ix3218 (.Y (nx3217), .A0 (nx4119), .A1 (nx7785), .B0 (nx4124)) ;
    nor03_2x ix4120 (.Y (nx4119), .A0 (nx396), .A1 (nx7427), .A2 (nx7401)) ;
    nand02 ix375 (.Y (nx374), .A0 (nx3925), .A1 (CNNIMGLOAD)) ;
    nand04 ix4125 (.Y (nx4124), .A0 (i8_counterout2_1), .A1 (nx7811), .A2 (
           nx7395), .A3 (nx7777)) ;
    nand03 ix423 (.Y (nx3102), .A0 (nx3940), .A1 (nx4126), .A2 (nx7961)) ;
    inv01 ix3238 (.Y (nx3237), .A (nx4131)) ;
    nor02_2x ix4132 (.Y (nx4131), .A0 (nx3233), .A1 (nx3235)) ;
    nor02_2x ix3234 (.Y (nx3233), .A0 (nx7815), .A1 (nx7419)) ;
    dff reg_i8_counterout2_3 (.Q (i8_counterout2_3), .QB (\$dummy [5]), .D (
        nx3237), .CLK (CLK)) ;
    aoi32 ix3236 (.Y (nx3235), .A0 (nx7811), .A1 (nx7395), .A2 (nx7777), .B0 (
          nx4138), .B1 (nx3101)) ;
    nor03_2x ix4139 (.Y (nx4138), .A0 (nx424), .A1 (nx7427), .A2 (nx7401)) ;
    nor02_2x ix425 (.Y (nx424), .A0 (nx7815), .A1 (nx4141)) ;
    nor03_2x ix4142 (.Y (nx4141), .A0 (i8_counterout2_0), .A1 (i8_counterout2_1)
             , .A2 (nx7911)) ;
    nand03 ix439 (.Y (nx3101), .A0 (nx7813), .A1 (nx7961), .A2 (nx7815)) ;
    dff reg_i8_counterout2_4 (.Q (i8_counterout2_4), .QB (nx4151), .D (nx3247), 
        .CLK (CLK)) ;
    inv01 ix3248 (.Y (nx3247), .A (nx4148)) ;
    aoi44 ix4149 (.Y (nx4148), .A0 (i8_counterout2_4), .A1 (nx7811), .A2 (nx7395
          ), .A3 (nx7777), .B0 (nx3947), .B1 (nx7737), .B2 (nx444), .B3 (nx7419)
          ) ;
    nand03 ix515 (.Y (nx514), .A0 (i8_counterout2_6), .A1 (i8_counterout2_7), .A2 (
           i8_counterout2_5)) ;
    dff reg_i8_counterout2_6 (.Q (i8_counterout2_6), .QB (nx4167), .D (nx3267), 
        .CLK (CLK)) ;
    inv01 ix3268 (.Y (nx3267), .A (nx4155)) ;
    aoi44 ix4156 (.Y (nx4155), .A0 (i8_counterout2_6), .A1 (nx7811), .A2 (nx7395
          ), .A3 (nx7777), .B0 (nx3947), .B1 (nx7737), .B2 (nx480), .B3 (nx7419)
          ) ;
    nand04 ix459 (.Y (nx458), .A0 (nx4141), .A1 (nx7815), .A2 (nx4151), .A3 (
           nx4159)) ;
    inv01 ix3258 (.Y (nx3257), .A (nx4162)) ;
    aoi44 ix4163 (.Y (nx4162), .A0 (i8_counterout2_5), .A1 (nx4107), .A2 (nx7397
          ), .A3 (nx7777), .B0 (nx3947), .B1 (nx7737), .B2 (nx464), .B3 (nx7419)
          ) ;
    dff reg_i8_counterout2_5 (.Q (i8_counterout2_5), .QB (nx4159), .D (nx3257), 
        .CLK (CLK)) ;
    nand04 ix457 (.Y (nx3100), .A0 (nx7813), .A1 (nx7961), .A2 (nx7815), .A3 (
           nx4151)) ;
    dff reg_i8_counterout2_7 (.Q (i8_counterout2_7), .QB (nx4177), .D (nx3277), 
        .CLK (CLK)) ;
    inv01 ix3278 (.Y (nx3277), .A (nx4171)) ;
    aoi44 ix4172 (.Y (nx4171), .A0 (i8_counterout2_7), .A1 (nx4107), .A2 (nx7397
          ), .A3 (nx7779), .B0 (nx494), .B1 (nx3947), .B2 (nx7739), .B3 (nx7419)
          ) ;
    nand04 ix4180 (.Y (nx4179), .A0 (i8_counterout2_0), .A1 (nx7811), .A2 (
           nx7397), .A3 (nx7779)) ;
    nor03_2x ix4182 (.Y (nx4181), .A0 (nx4167), .A1 (nx4177), .A2 (nx4159)) ;
    nor02_2x ix589 (.Y (nx588), .A0 (i8_loadenableD), .A1 (nx3917)) ;
    dff i8_reg_loadenableD (.Q (i8_loadenableD), .QB (\$dummy [6]), .D (
        loadingCNN), .CLK (CLK)) ;
    nand02 ix4189 (.Y (nx4188), .A0 (nx4191), .A1 (nx7415)) ;
    inv01 ix4192 (.Y (nx4191), .A (DataBus[14])) ;
    nor03_2x ix129 (.Y (nx128), .A0 (i8_counterout1_0), .A1 (nx102), .A2 (nx7401
             )) ;
    nand02 ix103 (.Y (nx102), .A0 (nx7771), .A1 (CNNIMGLOAD)) ;
    oai21 ix4197 (.Y (nx4196), .A0 (nx3917), .A1 (nx4029), .B0 (i8_counterout1_0
          )) ;
    oai21 ix603 (.Y (nx602), .A0 (zed), .A1 (nx362), .B0 (nx54)) ;
    nor02_2x ix3484 (.Y (nx3483), .A0 (nx4203), .A1 (nx1154)) ;
    dffs_ni i7_reg_read1 (.Q (EnableReadingFromCPU1), .QB (nx4203), .D (nx3483)
            , .CLK (CLK), .S (nx1158)) ;
    nand02 ix1159 (.Y (nx1158), .A0 (nx1154), .A1 (nx7823)) ;
    nand04 ix1155 (.Y (nx1154), .A0 (nx4207), .A1 (nx4370), .A2 (nx4447), .A3 (
           nx4277)) ;
    nor03_2x ix4208 (.Y (nx4207), .A0 (nx4209), .A1 (i7_counterout1_1), .A2 (
             nx1130)) ;
    oai21 ix3408 (.Y (nx3407), .A0 (nx4212), .A1 (nx7835), .B0 (nx4517)) ;
    nor02_2x ix4213 (.Y (nx4212), .A0 (nx960), .A1 (nx952)) ;
    oai21 ix961 (.Y (nx960), .A0 (nx4209), .A1 (nx4215), .B0 (nx4509)) ;
    oai21 ix4216 (.Y (nx4215), .A0 (CNNIMGLOAD), .A1 (nx7401), .B0 (nx4217)) ;
    nor03_2x ix639 (.Y (nx638), .A0 (CNNIMGLOAD), .A1 (nx7957), .A2 (nx4220)) ;
    nand02 ix4221 (.Y (nx4220), .A0 (nx7823), .A1 (nx4203)) ;
    nor02_2x ix3394 (.Y (nx3393), .A0 (nx7819), .A1 (nx836)) ;
    nor02_2x ix837 (.Y (nx836), .A0 (nx4217), .A1 (nx4227)) ;
    nor03_2x ix831 (.Y (nx830), .A0 (CNNIMGLOAD), .A1 (nx7957), .A2 (nx4231)) ;
    nand02 ix4232 (.Y (nx4231), .A0 (nx7819), .A1 (nx4233)) ;
    nor02_2x ix3384 (.Y (nx3383), .A0 (nx4233), .A1 (nx814)) ;
    nand04 ix815 (.Y (nx814), .A0 (nx4237), .A1 (nx4281), .A2 (nx4343), .A3 (
           nx4277)) ;
    nor03_2x ix4238 (.Y (nx4237), .A0 (nx4239), .A1 (nx4318), .A2 (nx802)) ;
    inv01 ix3328 (.Y (nx3327), .A (nx4243)) ;
    aoi44 ix4244 (.Y (nx4243), .A0 (i7_counterout2_2), .A1 (nx7827), .A2 (nx7392
          ), .A3 (nx7821), .B0 (nx4301), .B1 (nx7739), .B2 (nx690), .B3 (nx650)
          ) ;
    dff reg_i7_counterout2_2 (.Q (i7_counterout2_2), .QB (nx4239), .D (nx3327), 
        .CLK (CLK)) ;
    nand02 ix4247 (.Y (nx4246), .A0 (i7_reset2), .A1 (i7_tmp)) ;
    dffr i7_ix81 (.Q (i7_reset2), .QB (nx4227), .D (nx2), .CLK (CLK), .R (nx830)
         ) ;
    nor02_2x ix1141 (.Y (nx1140), .A0 (nx4251), .A1 (nx4501)) ;
    nor03_2x ix4252 (.Y (nx4251), .A0 (nx1134), .A1 (nx1130), .A2 (nx1128)) ;
    nand02 ix1135 (.Y (nx1134), .A0 (i7_counterout1_0), .A1 (nx4255)) ;
    dff reg_i7_counterout1_0 (.Q (i7_counterout1_0), .QB (nx4209), .D (nx3407), 
        .CLK (CLK)) ;
    oai21 ix3418 (.Y (nx3417), .A0 (nx4258), .A1 (nx7833), .B0 (nx4496)) ;
    aoi322 ix4259 (.Y (nx4258), .A0 (nx940), .A1 (nx4263), .A2 (nx7441), .B0 (
           nx4267), .B1 (nx7829), .C0 (i7_counterout1_1), .C1 (nx974)) ;
    inv01 ix941 (.Y (nx940), .A (nx4261)) ;
    nor02_2x ix4262 (.Y (nx4261), .A0 (DataBus[9]), .A1 (DataBus[8])) ;
    nand02 ix4264 (.Y (nx4263), .A0 (DataBus[8]), .A1 (DataBus[9])) ;
    dffr i7_ix59 (.Q (\$dummy [7]), .QB (nx4217), .D (nx2), .CLK (CLK), .R (
         nx638)) ;
    nor02_2x ix4268 (.Y (nx4267), .A0 (i7_counterout1_0), .A1 (i7_counterout1_1)
             ) ;
    dff reg_i7_counterout1_1 (.Q (i7_counterout1_1), .QB (nx4255), .D (nx3417), 
        .CLK (CLK)) ;
    nor03_2x ix4272 (.Y (nx4271), .A0 (nx7441), .A1 (CNNIMGLOAD), .A2 (nx7403)
             ) ;
    mux21 ix975 (.Y (nx974), .A0 (nx7441), .A1 (nx4209), .S0 (nx7829)) ;
    oai21 ix4275 (.Y (nx4274), .A0 (nx856), .A1 (i7_start), .B0 (loadingimg)) ;
    oai21 ix857 (.Y (nx856), .A0 (nx4217), .A1 (nx4277), .B0 (i7_read2)) ;
    nor03_2x ix1149 (.Y (nx1148), .A0 (nx812), .A1 (nx4367), .A2 (nx1138)) ;
    nand03 ix813 (.Y (nx812), .A0 (nx4237), .A1 (nx4281), .A2 (nx4343)) ;
    nor02_2x ix4282 (.Y (nx4281), .A0 (nx4283), .A1 (nx4333)) ;
    oai21 ix3348 (.Y (nx3347), .A0 (nx4287), .A1 (nx7839), .B0 (nx4331)) ;
    nor03_2x ix4288 (.Y (nx4287), .A0 (nx724), .A1 (nx7447), .A2 (nx7403)) ;
    dff reg_i7_counterout2_4 (.Q (i7_counterout2_4), .QB (nx4283), .D (nx3347), 
        .CLK (CLK)) ;
    nand03 ix719 (.Y (nx3111), .A0 (nx7837), .A1 (nx4239), .A2 (nx4318)) ;
    nor02_2x ix4294 (.Y (nx4293), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)
             ) ;
    dff reg_i7_counterout2_0 (.Q (i7_counterout2_0), .QB (nx4309), .D (nx3307), 
        .CLK (CLK)) ;
    oai21 ix3308 (.Y (nx3307), .A0 (nx4298), .A1 (nx7839), .B0 (nx4307)) ;
    nand02 ix655 (.Y (nx654), .A0 (nx4301), .A1 (nx7739)) ;
    nor02_2x ix4302 (.Y (nx4301), .A0 (i7_reset2), .A1 (CNNIMGLOAD)) ;
    oai21 ix649 (.Y (nx648), .A0 (nx4227), .A1 (nx4277), .B0 (nx7390)) ;
    nand04 ix4308 (.Y (nx4307), .A0 (i7_counterout2_0), .A1 (nx7825), .A2 (
           nx7390), .A3 (nx7819)) ;
    dff reg_i7_counterout2_1 (.Q (i7_counterout2_1), .QB (nx4317), .D (nx3317), 
        .CLK (CLK)) ;
    oai21 ix3318 (.Y (nx3317), .A0 (nx4312), .A1 (nx7839), .B0 (nx4315)) ;
    nor04 ix4313 (.Y (nx4312), .A0 (nx674), .A1 (i7_reset2), .A2 (CNNIMGLOAD), .A3 (
          nx7403)) ;
    nand04 ix4316 (.Y (nx4315), .A0 (i7_counterout2_1), .A1 (nx7825), .A2 (
           nx7390), .A3 (nx7819)) ;
    oai21 ix3338 (.Y (nx3337), .A0 (nx4322), .A1 (nx7839), .B0 (nx4327)) ;
    nor04 ix4323 (.Y (nx4322), .A0 (nx708), .A1 (i7_reset2), .A2 (CNNIMGLOAD), .A3 (
          nx7403)) ;
    dff reg_i7_counterout2_3 (.Q (i7_counterout2_3), .QB (nx4318), .D (nx3337), 
        .CLK (CLK)) ;
    nand04 ix4328 (.Y (nx4327), .A0 (i7_counterout2_3), .A1 (nx7825), .A2 (
           nx7390), .A3 (nx7819)) ;
    nand04 ix4332 (.Y (nx4331), .A0 (i7_counterout2_4), .A1 (nx7825), .A2 (
           nx7390), .A3 (nx7819)) ;
    inv01 ix3358 (.Y (nx3357), .A (nx4336)) ;
    aoi44 ix4337 (.Y (nx4336), .A0 (i7_counterout2_5), .A1 (nx7825), .A2 (nx7390
          ), .A3 (nx7821), .B0 (nx4301), .B1 (nx7739), .B2 (nx740), .B3 (nx650)
          ) ;
    dff reg_i7_counterout2_5 (.Q (i7_counterout2_5), .QB (nx4333), .D (nx3357), 
        .CLK (CLK)) ;
    nand04 ix735 (.Y (nx3109), .A0 (nx7837), .A1 (nx4239), .A2 (nx4318), .A3 (
           nx4283)) ;
    nand03 ix651 (.Y (nx650), .A0 (nx7825), .A1 (nx7390), .A2 (nx7821)) ;
    nor02_2x ix4344 (.Y (nx4343), .A0 (nx4345), .A1 (nx4355)) ;
    inv01 ix3368 (.Y (nx3367), .A (nx4348)) ;
    aoi44 ix4349 (.Y (nx4348), .A0 (i7_counterout2_6), .A1 (nx7825), .A2 (nx7392
          ), .A3 (nx7821), .B0 (nx4301), .B1 (nx7739), .B2 (nx758), .B3 (nx650)
          ) ;
    dff reg_i7_counterout2_6 (.Q (i7_counterout2_6), .QB (nx4345), .D (nx3367), 
        .CLK (CLK)) ;
    nand04 ix753 (.Y (nx3107), .A0 (nx4353), .A1 (nx4318), .A2 (nx4283), .A3 (
           nx4333)) ;
    nor03_2x ix4354 (.Y (nx4353), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)
             , .A2 (i7_counterout2_2)) ;
    inv01 ix3378 (.Y (nx3377), .A (nx4359)) ;
    aoi44 ix4360 (.Y (nx4359), .A0 (i7_counterout2_7), .A1 (nx7827), .A2 (nx7392
          ), .A3 (nx7821), .B0 (nx4301), .B1 (nx7739), .B2 (nx772), .B3 (nx650)
          ) ;
    dff reg_i7_counterout2_7 (.Q (i7_counterout2_7), .QB (nx4355), .D (nx3377), 
        .CLK (CLK)) ;
    nand02 ix4368 (.Y (nx4367), .A0 (nx7441), .A1 (i7_reset2)) ;
    nand03 ix1139 (.Y (nx1138), .A0 (nx4207), .A1 (nx4370), .A2 (nx4447)) ;
    nor02_2x ix4371 (.Y (nx4370), .A0 (i7_counterout1_4), .A1 (i7_counterout1_5)
             ) ;
    oai21 ix3448 (.Y (nx3447), .A0 (nx4374), .A1 (nx7833), .B0 (nx4430)) ;
    aoi322 ix4375 (.Y (nx4374), .A0 (nx894), .A1 (nx4383), .A2 (nx7441), .B0 (
           nx4386), .B1 (nx7829), .C0 (i7_counterout1_4), .C1 (nx1034)) ;
    oai21 ix895 (.Y (nx894), .A0 (nx4377), .A1 (nx4379), .B0 (nx4381)) ;
    inv02 ix4378 (.Y (nx4377), .A (DataBus[11])) ;
    nand03 ix4380 (.Y (nx4379), .A0 (DataBus[10]), .A1 (DataBus[8]), .A2 (
           DataBus[9])) ;
    inv02 ix4382 (.Y (nx4381), .A (DataBus[12])) ;
    nand03 ix1029 (.Y (nx3117), .A0 (nx4267), .A1 (nx4389), .A2 (nx4409)) ;
    oai21 ix3428 (.Y (nx3427), .A0 (nx4393), .A1 (nx7833), .B0 (nx4403)) ;
    aoi322 ix4394 (.Y (nx4393), .A0 (nx926), .A1 (nx4379), .A2 (nx7441), .B0 (
           nx4399), .B1 (nx7829), .C0 (i7_counterout1_2), .C1 (nx994)) ;
    nand02 ix927 (.Y (nx926), .A0 (nx4263), .A1 (nx4397)) ;
    inv01 ix4398 (.Y (nx4397), .A (DataBus[10])) ;
    nor03_2x ix4400 (.Y (nx4399), .A0 (i7_counterout1_0), .A1 (i7_counterout1_1)
             , .A2 (i7_counterout1_2)) ;
    dff reg_i7_counterout1_2 (.Q (i7_counterout1_2), .QB (nx4389), .D (nx3427), 
        .CLK (CLK)) ;
    mux21 ix995 (.Y (nx994), .A0 (nx7441), .A1 (nx4267), .S0 (nx7829)) ;
    oai21 ix4404 (.Y (nx4403), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_2
          )) ;
    nand02 ix4406 (.Y (nx4405), .A0 (nx7741), .A1 (nx7907)) ;
    oai21 ix3438 (.Y (nx3437), .A0 (nx4413), .A1 (nx7833), .B0 (nx4425)) ;
    aoi322 ix4414 (.Y (nx4413), .A0 (nx912), .A1 (nx4417), .A2 (nx7443), .B0 (
           nx4419), .B1 (nx7829), .C0 (i7_counterout1_3), .C1 (nx1014)) ;
    oai21 ix913 (.Y (nx912), .A0 (nx4397), .A1 (nx4263), .B0 (nx4377)) ;
    nand04 ix4418 (.Y (nx4417), .A0 (DataBus[11]), .A1 (DataBus[10]), .A2 (
           DataBus[8]), .A3 (DataBus[9])) ;
    nand03 ix1009 (.Y (nx3118), .A0 (nx4209), .A1 (nx4255), .A2 (nx4389)) ;
    dff reg_i7_counterout1_3 (.Q (i7_counterout1_3), .QB (nx4409), .D (nx3437), 
        .CLK (CLK)) ;
    mux21 ix1015 (.Y (nx1014), .A0 (nx7443), .A1 (nx4399), .S0 (nx7829)) ;
    oai21 ix4426 (.Y (nx4425), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_3
          )) ;
    dff reg_i7_counterout1_4 (.Q (i7_counterout1_4), .QB (nx4427), .D (nx3447), 
        .CLK (CLK)) ;
    mux21 ix1035 (.Y (nx1034), .A0 (nx7443), .A1 (nx4419), .S0 (nx7831)) ;
    oai21 ix4431 (.Y (nx4430), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_4
          )) ;
    oai21 ix3458 (.Y (nx3457), .A0 (nx4434), .A1 (nx7833), .B0 (nx4445)) ;
    aoi222 ix4435 (.Y (nx4434), .A0 (nx1058), .A1 (nx7443), .B0 (nx4437), .B1 (
           nx7831), .C0 (i7_counterout1_5), .C1 (nx1054)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (DataBus[13]), .A1 (nx4383)) ;
    nand04 ix1049 (.Y (nx3116), .A0 (nx4267), .A1 (nx4389), .A2 (nx4409), .A3 (
           nx4427)) ;
    dff reg_i7_counterout1_5 (.Q (i7_counterout1_5), .QB (nx4441), .D (nx3457), 
        .CLK (CLK)) ;
    mux21 ix1055 (.Y (nx1054), .A0 (nx7443), .A1 (nx4386), .S0 (nx7831)) ;
    oai21 ix4446 (.Y (nx4445), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_5
          )) ;
    nor02_2x ix4448 (.Y (nx4447), .A0 (i7_counterout1_6), .A1 (i7_counterout1_7)
             ) ;
    oai21 ix3468 (.Y (nx3467), .A0 (nx4453), .A1 (nx7833), .B0 (nx4469)) ;
    aoi222 ix4454 (.Y (nx4453), .A0 (nx1084), .A1 (nx7443), .B0 (nx4462), .B1 (
           nx7831), .C0 (i7_counterout1_6), .C1 (nx1078)) ;
    inv01 ix1085 (.Y (nx1084), .A (nx4457)) ;
    xnor2 ix4458 (.Y (nx4457), .A0 (DataBus[14]), .A1 (nx1082)) ;
    nor03_2x ix1083 (.Y (nx1082), .A0 (nx4460), .A1 (nx4381), .A2 (nx4417)) ;
    inv01 ix4461 (.Y (nx4460), .A (DataBus[13])) ;
    nand04 ix1073 (.Y (nx3115), .A0 (nx4399), .A1 (nx4409), .A2 (nx4427), .A3 (
           nx4441)) ;
    dff reg_i7_counterout1_6 (.Q (i7_counterout1_6), .QB (nx4465), .D (nx3467), 
        .CLK (CLK)) ;
    mux21 ix1079 (.Y (nx1078), .A0 (nx7443), .A1 (nx4437), .S0 (nx7831)) ;
    oai21 ix4470 (.Y (nx4469), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_6
          )) ;
    dff reg_i7_counterout1_7 (.Q (i7_counterout1_7), .QB (nx4487), .D (nx3477), 
        .CLK (CLK)) ;
    oai21 ix3478 (.Y (nx3477), .A0 (nx4475), .A1 (nx7833), .B0 (nx4485)) ;
    aoi222 ix4476 (.Y (nx4475), .A0 (nx1110), .A1 (nx7445), .B0 (nx1100), .B1 (
           nx7831), .C0 (i7_counterout1_7), .C1 (nx874)) ;
    xnor2 ix1111 (.Y (nx1110), .A0 (DataBus[15]), .A1 (nx4479)) ;
    nand02 ix4480 (.Y (nx4479), .A0 (DataBus[14]), .A1 (nx1082)) ;
    nor02_2x ix875 (.Y (nx874), .A0 (nx7445), .A1 (nx7831)) ;
    oai21 ix4486 (.Y (nx4485), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_7
          )) ;
    dffs_ni i7_reg_read2 (.Q (i7_read2), .QB (nx4233), .D (nx3383), .CLK (CLK), 
            .S (nx818)) ;
    nand02 ix819 (.Y (nx818), .A0 (nx814), .A1 (nx7821)) ;
    dffs_ni i7_reg_start (.Q (i7_start), .QB (\$dummy [8]), .D (nx3393), .CLK (
            CLK), .S (nx846)) ;
    nor03_2x ix847 (.Y (nx846), .A0 (i7_loadenableD), .A1 (CNNIMGLOAD), .A2 (
             nx7957)) ;
    dff i7_reg_loadenableD (.Q (i7_loadenableD), .QB (\$dummy [9]), .D (
        loadingimg), .CLK (CLK)) ;
    oai21 ix4497 (.Y (nx4496), .A0 (nx7843), .A1 (nx7847), .B0 (i7_counterout1_1
          )) ;
    nand02 ix1131 (.Y (nx1130), .A0 (nx4389), .A1 (nx4409)) ;
    nand03 ix1129 (.Y (nx1128), .A0 (nx4370), .A1 (nx4465), .A2 (nx4487)) ;
    nor03_2x ix4502 (.Y (nx4501), .A0 (nx808), .A1 (nx802), .A2 (nx796)) ;
    nand02 ix809 (.Y (nx808), .A0 (i7_counterout2_2), .A1 (i7_counterout2_3)) ;
    nand02 ix803 (.Y (nx802), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)) ;
    nand03 ix797 (.Y (nx796), .A0 (nx4281), .A1 (i7_counterout2_6), .A2 (
           i7_counterout2_7)) ;
    nand02 ix4510 (.Y (nx4509), .A0 (nx4511), .A1 (nx7445)) ;
    inv01 ix4512 (.Y (nx4511), .A (DataBus[8])) ;
    nor03_2x ix953 (.Y (nx952), .A0 (i7_counterout1_0), .A1 (nx862), .A2 (nx7403
             )) ;
    nand02 ix863 (.Y (nx862), .A0 (nx4217), .A1 (nx7741)) ;
    oai21 ix4518 (.Y (nx4517), .A0 (nx7845), .A1 (nx7849), .B0 (i7_counterout1_0
          )) ;
    nor02ii ix2123 (.Y (nx2122), .A0 (nx7537), .A1 (nx7455)) ;
    nand02 ix2109 (.Y (nx2108), .A0 (nx4522), .A1 (nx7853)) ;
    nand04 ix4523 (.Y (nx4522), .A0 (nx4525), .A1 (nx7765), .A2 (nx7435), .A3 (
           nx7813)) ;
    nor02_2x ix4526 (.Y (nx4525), .A0 (nx7911), .A1 (i8_counterout2_3)) ;
    nor02_2x ix1189 (.Y (nx1188), .A0 (nx4532), .A1 (nx7785)) ;
    inv01 ix4533 (.Y (nx4532), .A (DataBus[0])) ;
    nand02 ix2119 (.Y (nx2118), .A0 (nx4535), .A1 (nx4537)) ;
    nand03 ix4536 (.Y (nx4535), .A0 (nx7813), .A1 (nx7419), .A2 (nx4525)) ;
    nor03_2x ix4538 (.Y (nx4537), .A0 (nx2106), .A1 (nx7427), .A2 (nx7403)) ;
    nor02_2x ix2107 (.Y (nx2106), .A0 (nx2098), .A1 (nx4542)) ;
    nand02 ix2099 (.Y (nx2098), .A0 (nx7961), .A1 (nx7815)) ;
    nand03 ix4543 (.Y (nx4542), .A0 (nx7765), .A1 (nx7435), .A2 (nx7813)) ;
    nor02ii ix2149 (.Y (nx2148), .A0 (nx7537), .A1 (nx7459)) ;
    nor02_2x ix1203 (.Y (nx1202), .A0 (nx4547), .A1 (nx7785)) ;
    inv01 ix4548 (.Y (nx4547), .A (DataBus[1])) ;
    nor02ii ix2175 (.Y (nx2174), .A0 (nx7537), .A1 (nx7463)) ;
    nor02_2x ix1217 (.Y (nx1216), .A0 (nx4553), .A1 (nx7785)) ;
    inv01 ix4554 (.Y (nx4553), .A (DataBus[2])) ;
    nor02ii ix2201 (.Y (nx2200), .A0 (nx7537), .A1 (nx7467)) ;
    nor02_2x ix1231 (.Y (nx1230), .A0 (nx4558), .A1 (nx7785)) ;
    inv01 ix4559 (.Y (nx4558), .A (DataBus[3])) ;
    nor02ii ix2227 (.Y (nx2226), .A0 (nx7537), .A1 (nx7471)) ;
    nor02_2x ix1245 (.Y (nx1244), .A0 (nx4565), .A1 (nx7785)) ;
    inv01 ix4566 (.Y (nx4565), .A (DataBus[4])) ;
    nor02ii ix2253 (.Y (nx2252), .A0 (nx7537), .A1 (nx7475)) ;
    nor02_2x ix1259 (.Y (nx1258), .A0 (nx4570), .A1 (nx7787)) ;
    inv01 ix4571 (.Y (nx4570), .A (DataBus[5])) ;
    nor02ii ix2279 (.Y (nx2278), .A0 (nx7537), .A1 (nx7479)) ;
    nor02_2x ix1273 (.Y (nx1272), .A0 (nx4577), .A1 (nx7787)) ;
    inv01 ix4578 (.Y (nx4577), .A (DataBus[6])) ;
    nor02ii ix2305 (.Y (nx2304), .A0 (nx2108), .A1 (nx7483)) ;
    nor02_2x ix1287 (.Y (nx1286), .A0 (nx4582), .A1 (nx7787)) ;
    inv01 ix4583 (.Y (nx4582), .A (DataBus[7])) ;
    nor02ii ix2335 (.Y (nx2334), .A0 (nx2108), .A1 (nx7487)) ;
    nor02_2x ix1301 (.Y (nx1300), .A0 (nx4511), .A1 (nx7787)) ;
    nor02ii ix2359 (.Y (nx2358), .A0 (nx2108), .A1 (nx7491)) ;
    nor02_2x ix1315 (.Y (nx1314), .A0 (nx4592), .A1 (nx7787)) ;
    inv01 ix4593 (.Y (nx4592), .A (DataBus[9])) ;
    nor02ii ix2383 (.Y (nx2382), .A0 (nx2108), .A1 (nx7495)) ;
    nor02_2x ix1329 (.Y (nx1328), .A0 (nx4397), .A1 (nx7787)) ;
    nor02ii ix2407 (.Y (nx2406), .A0 (nx2108), .A1 (nx7499)) ;
    nor02_2x ix1343 (.Y (nx1342), .A0 (nx4377), .A1 (nx7787)) ;
    nor02ii ix2431 (.Y (nx2430), .A0 (nx2108), .A1 (nx7503)) ;
    nor02_2x ix1357 (.Y (nx1356), .A0 (nx4381), .A1 (nx7789)) ;
    latch i8_r1_lat_q_13 (.Q (DecompressedData2[15]), .D (nx2444), .CLK (nx7541)
          ) ;
    nor02ii ix2445 (.Y (nx2444), .A0 (nx2108), .A1 (nx7507)) ;
    nor02_2x ix1371 (.Y (nx1370), .A0 (nx4460), .A1 (nx7789)) ;
    nor02ii ix2525 (.Y (nx2524), .A0 (nx7575), .A1 (nx7455)) ;
    nand02 ix2515 (.Y (nx2514), .A0 (nx4613), .A1 (nx7853)) ;
    nand04 ix4614 (.Y (nx4613), .A0 (nx4525), .A1 (nx7765), .A2 (nx7435), .A3 (
           nx7863)) ;
    nor02_2x ix4616 (.Y (nx4615), .A0 (nx3940), .A1 (i8_counterout2_1)) ;
    nand02 ix2521 (.Y (nx2520), .A0 (nx4618), .A1 (nx4621)) ;
    nand03 ix4619 (.Y (nx4618), .A0 (nx7863), .A1 (nx7421), .A2 (nx4525)) ;
    nor03_2x ix4622 (.Y (nx4621), .A0 (nx2512), .A1 (nx7427), .A2 (nx7405)) ;
    nor02_2x ix2513 (.Y (nx2512), .A0 (nx2098), .A1 (nx4625)) ;
    nand03 ix4626 (.Y (nx4625), .A0 (nx7765), .A1 (nx7435), .A2 (nx7863)) ;
    nor02ii ix2549 (.Y (nx2548), .A0 (nx7575), .A1 (nx7459)) ;
    nor02ii ix2573 (.Y (nx2572), .A0 (nx7575), .A1 (nx7463)) ;
    nor02ii ix2597 (.Y (nx2596), .A0 (nx7575), .A1 (nx7467)) ;
    nor02ii ix2621 (.Y (nx2620), .A0 (nx7575), .A1 (nx7471)) ;
    nor02ii ix2645 (.Y (nx2644), .A0 (nx7575), .A1 (nx7475)) ;
    nor02ii ix2669 (.Y (nx2668), .A0 (nx7575), .A1 (nx7479)) ;
    nor02ii ix2693 (.Y (nx2692), .A0 (nx2514), .A1 (nx7483)) ;
    nor02ii ix2723 (.Y (nx2722), .A0 (nx2514), .A1 (nx7487)) ;
    nor02ii ix2747 (.Y (nx2746), .A0 (nx2514), .A1 (nx7491)) ;
    nor02ii ix2771 (.Y (nx2770), .A0 (nx2514), .A1 (nx7495)) ;
    nor02ii ix2795 (.Y (nx2794), .A0 (nx2514), .A1 (nx7499)) ;
    nor02ii ix2819 (.Y (nx2818), .A0 (nx2514), .A1 (nx7503)) ;
    latch i8_r2_lat_q_13 (.Q (DecompressedData2[31]), .D (nx2832), .CLK (nx7579)
          ) ;
    nor02ii ix2833 (.Y (nx2832), .A0 (nx2514), .A1 (nx7507)) ;
    nor02ii ix2915 (.Y (nx2914), .A0 (nx7587), .A1 (nx7455)) ;
    nand02 ix2905 (.Y (nx2904), .A0 (nx4663), .A1 (nx7853)) ;
    nand04 ix4664 (.Y (nx4663), .A0 (nx4525), .A1 (nx7765), .A2 (nx7435), .A3 (
           nx7865)) ;
    nor02_2x ix4666 (.Y (nx4665), .A0 (i8_counterout2_0), .A1 (nx4126)) ;
    nand02 ix2911 (.Y (nx2910), .A0 (nx4668), .A1 (nx4670)) ;
    nand03 ix4669 (.Y (nx4668), .A0 (nx7865), .A1 (nx7421), .A2 (nx4525)) ;
    nor03_2x ix4671 (.Y (nx4670), .A0 (nx2902), .A1 (nx7427), .A2 (nx7405)) ;
    nor02_2x ix2903 (.Y (nx2902), .A0 (nx2098), .A1 (nx4673)) ;
    nand03 ix4674 (.Y (nx4673), .A0 (nx7765), .A1 (nx7435), .A2 (nx7865)) ;
    nor02ii ix2939 (.Y (nx2938), .A0 (nx7587), .A1 (nx7459)) ;
    nor02ii ix2963 (.Y (nx2962), .A0 (nx7587), .A1 (nx7463)) ;
    nor02ii ix2987 (.Y (nx2986), .A0 (nx7587), .A1 (nx7467)) ;
    nor02ii ix3011 (.Y (nx3010), .A0 (nx7587), .A1 (nx7471)) ;
    nor02ii ix3035 (.Y (nx3034), .A0 (nx7587), .A1 (nx7475)) ;
    nor02ii ix3059 (.Y (nx3058), .A0 (nx7587), .A1 (nx7479)) ;
    nor02ii ix3083 (.Y (nx3082), .A0 (nx2904), .A1 (nx7483)) ;
    nor02ii ix3113 (.Y (nx3112), .A0 (nx2904), .A1 (nx7487)) ;
    nor02ii ix3137 (.Y (nx3136), .A0 (nx2904), .A1 (nx7491)) ;
    nor02ii ix3161 (.Y (nx3160), .A0 (nx2904), .A1 (nx7495)) ;
    nor02ii ix3185 (.Y (nx3184), .A0 (nx2904), .A1 (nx7499)) ;
    nor02ii ix3209 (.Y (nx3208), .A0 (nx2904), .A1 (nx7503)) ;
    latch i8_r3_lat_q_13 (.Q (DecompressedData2[47]), .D (nx3222), .CLK (nx7591)
          ) ;
    nor02ii ix3223 (.Y (nx3222), .A0 (nx2904), .A1 (nx7507)) ;
    nor02ii ix3303 (.Y (nx3302), .A0 (nx7599), .A1 (nx7455)) ;
    nand02 ix3293 (.Y (nx3292), .A0 (nx4711), .A1 (nx7853)) ;
    nand04 ix4712 (.Y (nx4711), .A0 (nx4525), .A1 (nx7767), .A2 (nx7435), .A3 (
           nx7781)) ;
    nand02 ix3299 (.Y (nx3298), .A0 (nx4715), .A1 (nx4717)) ;
    nand03 ix4716 (.Y (nx4715), .A0 (nx7781), .A1 (nx7421), .A2 (nx4525)) ;
    nor03_2x ix4718 (.Y (nx4717), .A0 (nx3290), .A1 (nx7427), .A2 (nx7405)) ;
    nor02_2x ix3291 (.Y (nx3290), .A0 (nx2098), .A1 (nx4720)) ;
    nand03 ix4721 (.Y (nx4720), .A0 (nx7767), .A1 (nx7437), .A2 (nx7781)) ;
    nor02ii ix3327 (.Y (nx3326), .A0 (nx7599), .A1 (nx7459)) ;
    nor02ii ix3351 (.Y (nx3350), .A0 (nx7599), .A1 (nx7463)) ;
    nor02ii ix3375 (.Y (nx3374), .A0 (nx7599), .A1 (nx7467)) ;
    nor02ii ix3399 (.Y (nx3398), .A0 (nx7599), .A1 (nx7471)) ;
    nor02ii ix3423 (.Y (nx3422), .A0 (nx7599), .A1 (nx7475)) ;
    nor02ii ix3447 (.Y (nx3446), .A0 (nx7599), .A1 (nx7479)) ;
    nor02ii ix3471 (.Y (nx3470), .A0 (nx3292), .A1 (nx7483)) ;
    nor02ii ix3501 (.Y (nx3500), .A0 (nx3292), .A1 (nx7487)) ;
    nor02ii ix3525 (.Y (nx3524), .A0 (nx3292), .A1 (nx7491)) ;
    nor02ii ix3549 (.Y (nx3548), .A0 (nx3292), .A1 (nx7495)) ;
    nor02ii ix3573 (.Y (nx3572), .A0 (nx3292), .A1 (nx7499)) ;
    nor02ii ix3597 (.Y (nx3596), .A0 (nx3292), .A1 (nx7503)) ;
    latch i8_r4_lat_q_13 (.Q (DecompressedData2[63]), .D (nx3610), .CLK (nx7603)
          ) ;
    nor02ii ix3611 (.Y (nx3610), .A0 (nx3292), .A1 (nx7507)) ;
    nor02ii ix3703 (.Y (nx3702), .A0 (nx7611), .A1 (nx7455)) ;
    nand02 ix3689 (.Y (nx3688), .A0 (nx4757), .A1 (nx7853)) ;
    nand04 ix4758 (.Y (nx4757), .A0 (nx4759), .A1 (nx7767), .A2 (nx7437), .A3 (
           nx7813)) ;
    nor02_2x ix4760 (.Y (nx4759), .A0 (nx7961), .A1 (i8_counterout2_3)) ;
    nand02 ix3699 (.Y (nx3698), .A0 (nx4763), .A1 (nx4765)) ;
    nand03 ix4764 (.Y (nx4763), .A0 (nx4114), .A1 (nx7421), .A2 (nx4759)) ;
    nor03_2x ix4766 (.Y (nx4765), .A0 (nx3686), .A1 (nx7429), .A2 (nx7405)) ;
    nor02_2x ix3687 (.Y (nx3686), .A0 (nx3682), .A1 (nx4542)) ;
    nand02 ix3683 (.Y (nx3682), .A0 (nx7911), .A1 (nx7815)) ;
    nor02ii ix3727 (.Y (nx3726), .A0 (nx7611), .A1 (nx7459)) ;
    nor02ii ix3751 (.Y (nx3750), .A0 (nx7611), .A1 (nx7463)) ;
    nor02ii ix3775 (.Y (nx3774), .A0 (nx7611), .A1 (nx7467)) ;
    nor02ii ix3799 (.Y (nx3798), .A0 (nx7611), .A1 (nx7471)) ;
    nor02ii ix3823 (.Y (nx3822), .A0 (nx7611), .A1 (nx7475)) ;
    nor02ii ix3847 (.Y (nx3846), .A0 (nx7611), .A1 (nx7479)) ;
    nor02ii ix3871 (.Y (nx3870), .A0 (nx3688), .A1 (nx7483)) ;
    nor02ii ix3901 (.Y (nx3900), .A0 (nx3688), .A1 (nx7487)) ;
    nor02ii ix3925 (.Y (nx3924), .A0 (nx3688), .A1 (nx7491)) ;
    nor02ii ix3949 (.Y (nx3948), .A0 (nx3688), .A1 (nx7495)) ;
    nor02ii ix3973 (.Y (nx3972), .A0 (nx3688), .A1 (nx7499)) ;
    nor02ii ix3997 (.Y (nx3996), .A0 (nx3688), .A1 (nx7503)) ;
    latch i8_r5_lat_q_13 (.Q (DecompressedData2[79]), .D (nx4010), .CLK (nx7615)
          ) ;
    nor02ii ix4011 (.Y (nx4010), .A0 (nx3688), .A1 (nx7507)) ;
    nor02ii ix4087 (.Y (nx4086), .A0 (nx7623), .A1 (nx7455)) ;
    nand02 ix4077 (.Y (nx4076), .A0 (nx4804), .A1 (nx7853)) ;
    nand04 ix4805 (.Y (nx4804), .A0 (nx4759), .A1 (nx7767), .A2 (nx7437), .A3 (
           nx7863)) ;
    nand02 ix4083 (.Y (nx4082), .A0 (nx4807), .A1 (nx4809)) ;
    nand03 ix4808 (.Y (nx4807), .A0 (nx7863), .A1 (nx7421), .A2 (nx4759)) ;
    nor03_2x ix4810 (.Y (nx4809), .A0 (nx4074), .A1 (nx7429), .A2 (nx7405)) ;
    nor02_2x ix4075 (.Y (nx4074), .A0 (nx3682), .A1 (nx4625)) ;
    nor02ii ix4111 (.Y (nx4110), .A0 (nx7623), .A1 (nx7459)) ;
    nor02ii ix4135 (.Y (nx4134), .A0 (nx7623), .A1 (nx7463)) ;
    nor02ii ix4159 (.Y (nx4158), .A0 (nx7623), .A1 (nx7467)) ;
    nor02ii ix4183 (.Y (nx4182), .A0 (nx7623), .A1 (nx7471)) ;
    nor02ii ix4207 (.Y (nx4206), .A0 (nx7623), .A1 (nx7475)) ;
    nor02ii ix4231 (.Y (nx4230), .A0 (nx7623), .A1 (nx7479)) ;
    nor02ii ix4255 (.Y (nx4254), .A0 (nx4076), .A1 (nx7483)) ;
    nor02ii ix4285 (.Y (nx4284), .A0 (nx4076), .A1 (nx7487)) ;
    nor02ii ix4309 (.Y (nx4308), .A0 (nx4076), .A1 (nx7491)) ;
    nor02ii ix4333 (.Y (nx4332), .A0 (nx4076), .A1 (nx7495)) ;
    nor02ii ix4357 (.Y (nx4356), .A0 (nx4076), .A1 (nx7499)) ;
    nor02ii ix4381 (.Y (nx4380), .A0 (nx4076), .A1 (nx7503)) ;
    latch i8_r6_lat_q_13 (.Q (DecompressedData2[95]), .D (nx4394), .CLK (nx7627)
          ) ;
    nor02ii ix4395 (.Y (nx4394), .A0 (nx4076), .A1 (nx7507)) ;
    nor02ii ix4481 (.Y (nx4480), .A0 (nx7643), .A1 (nx7455)) ;
    nand02 ix4471 (.Y (nx4470), .A0 (nx4847), .A1 (nx7853)) ;
    nand04 ix4848 (.Y (nx4847), .A0 (nx4759), .A1 (nx7767), .A2 (nx7437), .A3 (
           nx7865)) ;
    nand02 ix4477 (.Y (nx4476), .A0 (nx4851), .A1 (nx4853)) ;
    nand03 ix4852 (.Y (nx4851), .A0 (nx7865), .A1 (nx7421), .A2 (nx4759)) ;
    nor03_2x ix4854 (.Y (nx4853), .A0 (nx4468), .A1 (nx7429), .A2 (nx7405)) ;
    nor02_2x ix4469 (.Y (nx4468), .A0 (nx3682), .A1 (nx4673)) ;
    nor02ii ix4505 (.Y (nx4504), .A0 (nx7643), .A1 (nx7459)) ;
    nor02ii ix4529 (.Y (nx4528), .A0 (nx7643), .A1 (nx7463)) ;
    nor02ii ix4553 (.Y (nx4552), .A0 (nx7643), .A1 (nx7467)) ;
    nor02ii ix4577 (.Y (nx4576), .A0 (nx7643), .A1 (nx7471)) ;
    nor02ii ix4601 (.Y (nx4600), .A0 (nx7643), .A1 (nx7475)) ;
    nor02ii ix4625 (.Y (nx4624), .A0 (nx7643), .A1 (nx7479)) ;
    nor02ii ix4649 (.Y (nx4648), .A0 (nx4470), .A1 (nx7483)) ;
    nor02ii ix4679 (.Y (nx4678), .A0 (nx4470), .A1 (nx7487)) ;
    nor02ii ix4703 (.Y (nx4702), .A0 (nx4470), .A1 (nx7491)) ;
    nor02ii ix4727 (.Y (nx4726), .A0 (nx4470), .A1 (nx7495)) ;
    nor02ii ix4751 (.Y (nx4750), .A0 (nx4470), .A1 (nx7499)) ;
    nor02ii ix4775 (.Y (nx4774), .A0 (nx4470), .A1 (nx7503)) ;
    latch i8_r7_lat_q_13 (.Q (DecompressedData2[111]), .D (nx4788), .CLK (nx7647
          )) ;
    nor02ii ix4789 (.Y (nx4788), .A0 (nx4470), .A1 (nx7507)) ;
    nor02ii ix4865 (.Y (nx4864), .A0 (nx7655), .A1 (nx7457)) ;
    nand02 ix4855 (.Y (nx4854), .A0 (nx4894), .A1 (nx7855)) ;
    nand04 ix4895 (.Y (nx4894), .A0 (nx4759), .A1 (nx7767), .A2 (nx7437), .A3 (
           nx7781)) ;
    nand02 ix4861 (.Y (nx4860), .A0 (nx4897), .A1 (nx4899)) ;
    nand03 ix4898 (.Y (nx4897), .A0 (nx7781), .A1 (nx7421), .A2 (nx4759)) ;
    nor03_2x ix4900 (.Y (nx4899), .A0 (nx4852), .A1 (nx7429), .A2 (nx7405)) ;
    nor02_2x ix4853 (.Y (nx4852), .A0 (nx3682), .A1 (nx4720)) ;
    nor02ii ix4889 (.Y (nx4888), .A0 (nx7655), .A1 (nx7461)) ;
    nor02ii ix4913 (.Y (nx4912), .A0 (nx7655), .A1 (nx7465)) ;
    nor02ii ix4937 (.Y (nx4936), .A0 (nx7655), .A1 (nx7469)) ;
    nor02ii ix4961 (.Y (nx4960), .A0 (nx7655), .A1 (nx7473)) ;
    nor02ii ix4985 (.Y (nx4984), .A0 (nx7655), .A1 (nx7477)) ;
    nor02ii ix5009 (.Y (nx5008), .A0 (nx7655), .A1 (nx7481)) ;
    nor02ii ix5033 (.Y (nx5032), .A0 (nx4854), .A1 (nx7485)) ;
    nor02ii ix5063 (.Y (nx5062), .A0 (nx4854), .A1 (nx7489)) ;
    nor02ii ix5087 (.Y (nx5086), .A0 (nx4854), .A1 (nx7493)) ;
    nor02ii ix5111 (.Y (nx5110), .A0 (nx4854), .A1 (nx7497)) ;
    nor02ii ix5135 (.Y (nx5134), .A0 (nx4854), .A1 (nx7501)) ;
    nor02ii ix5159 (.Y (nx5158), .A0 (nx4854), .A1 (nx7505)) ;
    latch i8_r8_lat_q_13 (.Q (DecompressedData2[127]), .D (nx5172), .CLK (nx7659
          )) ;
    nor02ii ix5173 (.Y (nx5172), .A0 (nx4854), .A1 (nx7509)) ;
    nor02ii ix5263 (.Y (nx5262), .A0 (nx7667), .A1 (nx7457)) ;
    nand02 ix5249 (.Y (nx5248), .A0 (nx4937), .A1 (nx7855)) ;
    nand04 ix4938 (.Y (nx4937), .A0 (nx4939), .A1 (nx7767), .A2 (nx7437), .A3 (
           nx4114)) ;
    nor02_2x ix4940 (.Y (nx4939), .A0 (nx7911), .A1 (nx7817)) ;
    nand02 ix5259 (.Y (nx5258), .A0 (nx4942), .A1 (nx4945)) ;
    nand03 ix4943 (.Y (nx4942), .A0 (nx4114), .A1 (nx7423), .A2 (nx4939)) ;
    nor03_2x ix4946 (.Y (nx4945), .A0 (nx5246), .A1 (nx7429), .A2 (nx7407)) ;
    nor02_2x ix5247 (.Y (nx5246), .A0 (nx5242), .A1 (nx4542)) ;
    nand02 ix5243 (.Y (nx5242), .A0 (nx7809), .A1 (i8_counterout2_3)) ;
    nor02ii ix5287 (.Y (nx5286), .A0 (nx7667), .A1 (nx7461)) ;
    nor02ii ix5311 (.Y (nx5310), .A0 (nx7667), .A1 (nx7465)) ;
    nor02ii ix5335 (.Y (nx5334), .A0 (nx7667), .A1 (nx7469)) ;
    nor02ii ix5359 (.Y (nx5358), .A0 (nx7667), .A1 (nx7473)) ;
    nor02ii ix5383 (.Y (nx5382), .A0 (nx7667), .A1 (nx7477)) ;
    nor02ii ix5407 (.Y (nx5406), .A0 (nx7667), .A1 (nx7481)) ;
    nor02ii ix5431 (.Y (nx5430), .A0 (nx5248), .A1 (nx7485)) ;
    nor02ii ix5461 (.Y (nx5460), .A0 (nx5248), .A1 (nx7489)) ;
    nor02ii ix5485 (.Y (nx5484), .A0 (nx5248), .A1 (nx7493)) ;
    nor02ii ix5509 (.Y (nx5508), .A0 (nx5248), .A1 (nx7497)) ;
    nor02ii ix5533 (.Y (nx5532), .A0 (nx5248), .A1 (nx7501)) ;
    nor02ii ix5557 (.Y (nx5556), .A0 (nx5248), .A1 (nx7505)) ;
    latch i8_r9_lat_q_13 (.Q (DecompressedData2[143]), .D (nx5570), .CLK (nx7671
          )) ;
    nor02ii ix5571 (.Y (nx5570), .A0 (nx5248), .A1 (nx7509)) ;
    nor02ii ix5647 (.Y (nx5646), .A0 (nx7679), .A1 (nx7457)) ;
    nand02 ix5637 (.Y (nx5636), .A0 (nx4985), .A1 (nx7855)) ;
    nand04 ix4986 (.Y (nx4985), .A0 (nx4939), .A1 (nx3895), .A2 (nx7437), .A3 (
           nx7863)) ;
    nand02 ix5643 (.Y (nx5642), .A0 (nx4988), .A1 (nx4990)) ;
    nand03 ix4989 (.Y (nx4988), .A0 (nx7863), .A1 (nx7423), .A2 (nx4939)) ;
    nor03_2x ix4991 (.Y (nx4990), .A0 (nx5634), .A1 (nx7429), .A2 (nx7407)) ;
    nor02_2x ix5635 (.Y (nx5634), .A0 (nx5242), .A1 (nx4625)) ;
    nor02ii ix5671 (.Y (nx5670), .A0 (nx7679), .A1 (nx7461)) ;
    nor02ii ix5695 (.Y (nx5694), .A0 (nx7679), .A1 (nx7465)) ;
    nor02ii ix5719 (.Y (nx5718), .A0 (nx7679), .A1 (nx7469)) ;
    nor02ii ix5743 (.Y (nx5742), .A0 (nx7679), .A1 (nx7473)) ;
    nor02ii ix5767 (.Y (nx5766), .A0 (nx7679), .A1 (nx7477)) ;
    nor02ii ix5791 (.Y (nx5790), .A0 (nx7679), .A1 (nx7481)) ;
    nor02ii ix5815 (.Y (nx5814), .A0 (nx5636), .A1 (nx7485)) ;
    nor02ii ix5845 (.Y (nx5844), .A0 (nx5636), .A1 (nx7489)) ;
    nor02ii ix5869 (.Y (nx5868), .A0 (nx5636), .A1 (nx7493)) ;
    nor02ii ix5893 (.Y (nx5892), .A0 (nx5636), .A1 (nx7497)) ;
    nor02ii ix5917 (.Y (nx5916), .A0 (nx5636), .A1 (nx7501)) ;
    nor02ii ix5941 (.Y (nx5940), .A0 (nx5636), .A1 (nx7505)) ;
    latch i8_r10_lat_q_13 (.Q (DecompressedData2[159]), .D (nx5954), .CLK (
          nx7683)) ;
    nor02ii ix5955 (.Y (nx5954), .A0 (nx5636), .A1 (nx7509)) ;
    nor02ii ix6037 (.Y (nx6036), .A0 (nx7691), .A1 (nx7457)) ;
    nand02 ix6027 (.Y (nx6026), .A0 (nx5029), .A1 (nx7855)) ;
    nand04 ix5030 (.Y (nx5029), .A0 (nx4939), .A1 (nx3895), .A2 (nx7439), .A3 (
           nx7865)) ;
    nand02 ix6033 (.Y (nx6032), .A0 (nx5033), .A1 (nx5035)) ;
    nand03 ix5034 (.Y (nx5033), .A0 (nx7865), .A1 (nx7423), .A2 (nx4939)) ;
    nor03_2x ix5036 (.Y (nx5035), .A0 (nx6024), .A1 (nx7429), .A2 (nx7407)) ;
    nor02_2x ix6025 (.Y (nx6024), .A0 (nx5242), .A1 (nx4673)) ;
    nor02ii ix6061 (.Y (nx6060), .A0 (nx7691), .A1 (nx7461)) ;
    nor02ii ix6085 (.Y (nx6084), .A0 (nx7691), .A1 (nx7465)) ;
    nor02ii ix6109 (.Y (nx6108), .A0 (nx7691), .A1 (nx7469)) ;
    nor02ii ix6133 (.Y (nx6132), .A0 (nx7691), .A1 (nx7473)) ;
    nor02ii ix6157 (.Y (nx6156), .A0 (nx7691), .A1 (nx7477)) ;
    nor02ii ix6181 (.Y (nx6180), .A0 (nx7691), .A1 (nx7481)) ;
    nor02ii ix6205 (.Y (nx6204), .A0 (nx6026), .A1 (nx7485)) ;
    nor02ii ix6235 (.Y (nx6234), .A0 (nx6026), .A1 (nx7489)) ;
    nor02ii ix6259 (.Y (nx6258), .A0 (nx6026), .A1 (nx7493)) ;
    nor02ii ix6283 (.Y (nx6282), .A0 (nx6026), .A1 (nx7497)) ;
    nor02ii ix6307 (.Y (nx6306), .A0 (nx6026), .A1 (nx7501)) ;
    nor02ii ix6331 (.Y (nx6330), .A0 (nx6026), .A1 (nx7505)) ;
    latch i8_r11_lat_q_13 (.Q (DecompressedData2[175]), .D (nx6344), .CLK (
          nx7695)) ;
    nor02ii ix6345 (.Y (nx6344), .A0 (nx6026), .A1 (nx7509)) ;
    nor02ii ix6421 (.Y (nx6420), .A0 (nx7703), .A1 (nx7457)) ;
    nand02 ix6411 (.Y (nx6410), .A0 (nx5075), .A1 (nx7855)) ;
    nand04 ix5076 (.Y (nx5075), .A0 (nx4939), .A1 (nx3895), .A2 (nx7439), .A3 (
           nx3938)) ;
    nand02 ix6417 (.Y (nx6416), .A0 (nx5078), .A1 (nx5080)) ;
    nand03 ix5079 (.Y (nx5078), .A0 (nx3938), .A1 (nx7423), .A2 (nx4939)) ;
    nor03_2x ix5081 (.Y (nx5080), .A0 (nx6408), .A1 (nx7431), .A2 (nx7407)) ;
    nor02_2x ix6409 (.Y (nx6408), .A0 (nx5242), .A1 (nx4720)) ;
    nor02ii ix6445 (.Y (nx6444), .A0 (nx7703), .A1 (nx7461)) ;
    nor02ii ix6469 (.Y (nx6468), .A0 (nx7703), .A1 (nx7465)) ;
    nor02ii ix6493 (.Y (nx6492), .A0 (nx7703), .A1 (nx7469)) ;
    nor02ii ix6517 (.Y (nx6516), .A0 (nx7703), .A1 (nx7473)) ;
    nor02ii ix6541 (.Y (nx6540), .A0 (nx7703), .A1 (nx7477)) ;
    nor02ii ix6565 (.Y (nx6564), .A0 (nx7703), .A1 (nx7481)) ;
    nor02ii ix6589 (.Y (nx6588), .A0 (nx6410), .A1 (nx7485)) ;
    nor02ii ix6619 (.Y (nx6618), .A0 (nx6410), .A1 (nx7489)) ;
    nor02ii ix6643 (.Y (nx6642), .A0 (nx6410), .A1 (nx7493)) ;
    nor02ii ix6667 (.Y (nx6666), .A0 (nx6410), .A1 (nx7497)) ;
    nor02ii ix6691 (.Y (nx6690), .A0 (nx6410), .A1 (nx7501)) ;
    nor02ii ix6715 (.Y (nx6714), .A0 (nx6410), .A1 (nx7505)) ;
    latch i8_r12_lat_q_13 (.Q (DecompressedData2[191]), .D (nx6728), .CLK (
          nx7707)) ;
    nor02ii ix6729 (.Y (nx6728), .A0 (nx6410), .A1 (nx7509)) ;
    nor02ii ix6813 (.Y (nx6812), .A0 (nx7715), .A1 (nx7457)) ;
    nand02 ix6803 (.Y (nx6802), .A0 (nx5119), .A1 (nx7855)) ;
    nand04 ix5120 (.Y (nx5119), .A0 (nx5121), .A1 (nx3895), .A2 (nx7439), .A3 (
           nx4114)) ;
    nor02_2x ix5122 (.Y (nx5121), .A0 (nx7809), .A1 (nx7817)) ;
    nand02 ix6809 (.Y (nx6808), .A0 (nx5124), .A1 (nx5126)) ;
    nand03 ix5125 (.Y (nx5124), .A0 (nx4114), .A1 (nx5121), .A2 (nx7423)) ;
    nor03_2x ix5127 (.Y (nx5126), .A0 (nx6800), .A1 (nx7431), .A2 (nx7407)) ;
    nor02_2x ix6801 (.Y (nx6800), .A0 (nx520), .A1 (nx4542)) ;
    nand02 ix521 (.Y (nx520), .A0 (nx7911), .A1 (i8_counterout2_3)) ;
    nor02ii ix6837 (.Y (nx6836), .A0 (nx7715), .A1 (nx7461)) ;
    nor02ii ix6861 (.Y (nx6860), .A0 (nx7715), .A1 (nx7465)) ;
    nor02ii ix6885 (.Y (nx6884), .A0 (nx7715), .A1 (nx7469)) ;
    nor02ii ix6909 (.Y (nx6908), .A0 (nx7715), .A1 (nx7473)) ;
    nor02ii ix6933 (.Y (nx6932), .A0 (nx7715), .A1 (nx7477)) ;
    nor02ii ix6957 (.Y (nx6956), .A0 (nx7715), .A1 (nx7481)) ;
    nor02ii ix6981 (.Y (nx6980), .A0 (nx6802), .A1 (nx7485)) ;
    nor02ii ix7011 (.Y (nx7010), .A0 (nx6802), .A1 (nx7489)) ;
    nor02ii ix7035 (.Y (nx7034), .A0 (nx6802), .A1 (nx7493)) ;
    nor02ii ix7059 (.Y (nx7058), .A0 (nx6802), .A1 (nx7497)) ;
    nor02ii ix7083 (.Y (nx7082), .A0 (nx6802), .A1 (nx7501)) ;
    nor02ii ix7107 (.Y (nx7106), .A0 (nx6802), .A1 (nx7505)) ;
    latch i8_r13_lat_q_13 (.Q (DecompressedData2[207]), .D (nx7120), .CLK (
          nx7719)) ;
    nor02ii ix7121 (.Y (nx7120), .A0 (nx6802), .A1 (nx7509)) ;
    nor02ii ix7197 (.Y (nx7196), .A0 (nx7727), .A1 (nx7457)) ;
    nand02 ix7187 (.Y (nx7186), .A0 (nx5165), .A1 (nx7855)) ;
    nand04 ix5166 (.Y (nx5165), .A0 (nx5121), .A1 (nx3895), .A2 (nx7439), .A3 (
           nx4615)) ;
    nand02 ix7193 (.Y (nx7192), .A0 (nx5169), .A1 (nx5171)) ;
    nand03 ix5170 (.Y (nx5169), .A0 (nx4615), .A1 (nx5121), .A2 (nx7423)) ;
    nor03_2x ix5172 (.Y (nx5171), .A0 (nx7184), .A1 (nx7431), .A2 (nx7407)) ;
    nor02_2x ix7185 (.Y (nx7184), .A0 (nx520), .A1 (nx4625)) ;
    nor02ii ix7221 (.Y (nx7220), .A0 (nx7727), .A1 (nx7461)) ;
    nor02ii ix7245 (.Y (nx7244), .A0 (nx7727), .A1 (nx7465)) ;
    nor02ii ix7269 (.Y (nx7268), .A0 (nx7727), .A1 (nx7469)) ;
    nor02ii ix7293 (.Y (nx7292), .A0 (nx7727), .A1 (nx7473)) ;
    nor02ii ix7317 (.Y (nx7316), .A0 (nx7727), .A1 (nx7477)) ;
    nor02ii ix7341 (.Y (nx7340), .A0 (nx7727), .A1 (nx7481)) ;
    nor02ii ix7365 (.Y (nx7364), .A0 (nx7186), .A1 (nx7485)) ;
    nor02ii ix7395 (.Y (nx7394), .A0 (nx7186), .A1 (nx7489)) ;
    nor02ii ix7419 (.Y (nx7418), .A0 (nx7186), .A1 (nx7493)) ;
    nor02ii ix7443 (.Y (nx7442), .A0 (nx7186), .A1 (nx7497)) ;
    nor02ii ix7467 (.Y (nx7466), .A0 (nx7186), .A1 (nx7501)) ;
    nor02ii ix7491 (.Y (nx7490), .A0 (nx7186), .A1 (nx7505)) ;
    latch i8_r14_lat_q_13 (.Q (DecompressedData2[223]), .D (nx7504), .CLK (
          nx7731)) ;
    nor02ii ix7505 (.Y (nx7504), .A0 (nx7186), .A1 (nx7509)) ;
    nor02ii ix1193 (.Y (nx1192), .A0 (nx7451), .A1 (nx1188)) ;
    nand02 ix1177 (.Y (nx1176), .A0 (nx5209), .A1 (nx7857)) ;
    nand04 ix5210 (.Y (nx5209), .A0 (nx5121), .A1 (nx3895), .A2 (nx7439), .A3 (
           nx4665)) ;
    nand02 ix1187 (.Y (nx1186), .A0 (nx5212), .A1 (nx5215)) ;
    nand03 ix5213 (.Y (nx5212), .A0 (nx4665), .A1 (nx5121), .A2 (nx7423)) ;
    nor03_2x ix5216 (.Y (nx5215), .A0 (nx1174), .A1 (nx7431), .A2 (nx7407)) ;
    nor02_2x ix1175 (.Y (nx1174), .A0 (nx520), .A1 (nx4673)) ;
    nor02ii ix1207 (.Y (nx1206), .A0 (nx7451), .A1 (nx1202)) ;
    nor02ii ix1221 (.Y (nx1220), .A0 (nx7451), .A1 (nx1216)) ;
    nor02ii ix1235 (.Y (nx1234), .A0 (nx7451), .A1 (nx1230)) ;
    nor02ii ix1249 (.Y (nx1248), .A0 (nx7451), .A1 (nx1244)) ;
    nor02ii ix1263 (.Y (nx1262), .A0 (nx7451), .A1 (nx1258)) ;
    nor02ii ix1277 (.Y (nx1276), .A0 (nx7451), .A1 (nx1272)) ;
    nor02ii ix1291 (.Y (nx1290), .A0 (nx1176), .A1 (nx1286)) ;
    nor02ii ix1305 (.Y (nx1304), .A0 (nx1176), .A1 (nx1300)) ;
    nor02ii ix1319 (.Y (nx1318), .A0 (nx1176), .A1 (nx1314)) ;
    nor02ii ix1333 (.Y (nx1332), .A0 (nx1176), .A1 (nx1328)) ;
    nor02ii ix1347 (.Y (nx1346), .A0 (nx1176), .A1 (nx1342)) ;
    nor02ii ix1361 (.Y (nx1360), .A0 (nx1176), .A1 (nx1356)) ;
    nor02ii ix1375 (.Y (nx1374), .A0 (nx1176), .A1 (nx1370)) ;
    inv02 ix1389 (.Y (nx1388), .A (nx5259)) ;
    nor03_2x ix5260 (.Y (nx5259), .A0 (nx1386), .A1 (nx7431), .A2 (nx7409)) ;
    nor02ii ix1387 (.Y (nx1386), .A0 (nx4011), .A1 (nx5263)) ;
    nor03_2x ix5264 (.Y (nx5263), .A0 (nx3940), .A1 (nx4126), .A2 (nx520)) ;
    nand02 ix1395 (.Y (nx1394), .A0 (nx5266), .A1 (nx5259)) ;
    nand02 ix5267 (.Y (nx5266), .A0 (nx5263), .A1 (nx7425)) ;
    nor04 ix2087 (.Y (nx2086), .A0 (nx4532), .A1 (nx7839), .A2 (nx7447), .A3 (
          nx7409)) ;
    nand02 ix2081 (.Y (nx2080), .A0 (nx5303), .A1 (nx7869)) ;
    nand03 ix5304 (.Y (nx5303), .A0 (nx5305), .A1 (nx7529), .A2 (nx2072)) ;
    nor02_2x ix5306 (.Y (nx5305), .A0 (nx4309), .A1 (nx4317)) ;
    nor03_2x ix2069 (.Y (nx2068), .A0 (nx7845), .A1 (nx4283), .A2 (nx7839)) ;
    nor02_2x ix2073 (.Y (nx2072), .A0 (nx4318), .A1 (i7_counterout2_2)) ;
    nor04 ix2135 (.Y (nx2134), .A0 (nx4547), .A1 (nx7839), .A2 (nx7447), .A3 (
          nx7409)) ;
    nor04 ix2161 (.Y (nx2160), .A0 (nx4553), .A1 (nx7841), .A2 (nx7447), .A3 (
          nx7409)) ;
    nor04 ix2187 (.Y (nx2186), .A0 (nx4558), .A1 (nx7841), .A2 (nx7447), .A3 (
          nx7409)) ;
    nor04 ix2213 (.Y (nx2212), .A0 (nx4565), .A1 (nx7841), .A2 (nx7447), .A3 (
          nx7409)) ;
    nor04 ix2239 (.Y (nx2238), .A0 (nx4570), .A1 (nx7841), .A2 (nx7447), .A3 (
          nx7411)) ;
    nor04 ix2265 (.Y (nx2264), .A0 (nx4577), .A1 (nx7841), .A2 (nx7449), .A3 (
          nx7411)) ;
    nor04 ix2291 (.Y (nx2290), .A0 (nx4582), .A1 (nx7841), .A2 (nx7449), .A3 (
          nx7411)) ;
    nand02 ix2321 (.Y (nx2320), .A0 (nx5331), .A1 (nx7869)) ;
    nand03 ix5332 (.Y (nx5331), .A0 (nx5333), .A1 (nx7529), .A2 (nx2072)) ;
    nor02_2x ix5334 (.Y (nx5333), .A0 (i7_counterout2_0), .A1 (nx4317)) ;
    latch i7_r27_lat_q_5 (.Q (DecompressedData1[13]), .D (nx7553), .CLK (nx7571)
          ) ;
    latch i7_r27_lat_q_6 (.Q (DecompressedData1[14]), .D (nx7559), .CLK (nx7571)
          ) ;
    latch i7_r27_lat_q_7 (.Q (DecompressedData1[15]), .D (nx7565), .CLK (nx7571)
          ) ;
    nand02 ix2495 (.Y (nx2494), .A0 (nx5347), .A1 (nx7869)) ;
    nand03 ix5348 (.Y (nx5347), .A0 (nx5349), .A1 (nx7529), .A2 (nx2072)) ;
    nor02_2x ix5350 (.Y (nx5349), .A0 (nx4309), .A1 (i7_counterout2_1)) ;
    nand02 ix2709 (.Y (nx2708), .A0 (nx5362), .A1 (nx7869)) ;
    nand03 ix5363 (.Y (nx5362), .A0 (nx7837), .A1 (nx7529), .A2 (nx2072)) ;
    latch i7_r25_lat_q_5 (.Q (DecompressedData1[29]), .D (nx7553), .CLK (nx7583)
          ) ;
    latch i7_r25_lat_q_6 (.Q (DecompressedData1[30]), .D (nx7559), .CLK (nx7583)
          ) ;
    latch i7_r25_lat_q_7 (.Q (DecompressedData1[31]), .D (nx7565), .CLK (nx7583)
          ) ;
    nand02 ix2889 (.Y (nx2888), .A0 (nx5375), .A1 (nx7869)) ;
    nand03 ix5376 (.Y (nx5375), .A0 (nx5305), .A1 (nx7529), .A2 (nx2880)) ;
    nor02_2x ix2881 (.Y (nx2880), .A0 (i7_counterout2_3), .A1 (nx4239)) ;
    nand02 ix3099 (.Y (nx3098), .A0 (nx5389), .A1 (nx7869)) ;
    nand03 ix5390 (.Y (nx5389), .A0 (nx5333), .A1 (nx7529), .A2 (nx2880)) ;
    latch i7_r23_lat_q_5 (.Q (DecompressedData1[45]), .D (nx7553), .CLK (nx7595)
          ) ;
    latch i7_r23_lat_q_6 (.Q (DecompressedData1[46]), .D (nx7559), .CLK (nx7595)
          ) ;
    latch i7_r23_lat_q_7 (.Q (DecompressedData1[47]), .D (nx7565), .CLK (nx7595)
          ) ;
    nand02 ix3273 (.Y (nx3272), .A0 (nx5403), .A1 (nx7869)) ;
    nand03 ix5404 (.Y (nx5403), .A0 (nx5349), .A1 (nx7529), .A2 (nx2880)) ;
    nand02 ix3487 (.Y (nx3486), .A0 (nx5415), .A1 (nx7871)) ;
    nand03 ix5416 (.Y (nx5415), .A0 (nx7837), .A1 (nx7531), .A2 (nx2880)) ;
    latch i7_r21_lat_q_5 (.Q (DecompressedData1[61]), .D (nx7553), .CLK (nx7607)
          ) ;
    latch i7_r21_lat_q_6 (.Q (DecompressedData1[62]), .D (nx7559), .CLK (nx7607)
          ) ;
    latch i7_r21_lat_q_7 (.Q (DecompressedData1[63]), .D (nx7565), .CLK (nx7607)
          ) ;
    nand02 ix3669 (.Y (nx3668), .A0 (nx5427), .A1 (nx7871)) ;
    nand03 ix5428 (.Y (nx5427), .A0 (nx5305), .A1 (nx7531), .A2 (nx3660)) ;
    nor02_2x ix3661 (.Y (nx3660), .A0 (i7_counterout2_3), .A1 (i7_counterout2_2)
             ) ;
    nand02 ix3887 (.Y (nx3886), .A0 (nx5441), .A1 (nx7871)) ;
    nand03 ix5442 (.Y (nx5441), .A0 (nx5333), .A1 (nx7531), .A2 (nx3660)) ;
    latch i7_r19_lat_q_5 (.Q (DecompressedData1[77]), .D (nx7553), .CLK (nx7619)
          ) ;
    latch i7_r19_lat_q_6 (.Q (DecompressedData1[78]), .D (nx7559), .CLK (nx7619)
          ) ;
    latch i7_r19_lat_q_7 (.Q (DecompressedData1[79]), .D (nx7565), .CLK (nx7619)
          ) ;
    nand02 ix4061 (.Y (nx4060), .A0 (nx5454), .A1 (nx7871)) ;
    nand03 ix5455 (.Y (nx5454), .A0 (nx5349), .A1 (nx7531), .A2 (nx3660)) ;
    nand02 ix4271 (.Y (nx4270), .A0 (nx5467), .A1 (nx7871)) ;
    nand03 ix5468 (.Y (nx5467), .A0 (nx7837), .A1 (nx7531), .A2 (nx3660)) ;
    latch i7_r17_lat_q_5 (.Q (DecompressedData1[93]), .D (nx7553), .CLK (nx7631)
          ) ;
    latch i7_r17_lat_q_6 (.Q (DecompressedData1[94]), .D (nx7559), .CLK (nx7631)
          ) ;
    latch i7_r17_lat_q_7 (.Q (DecompressedData1[95]), .D (nx7565), .CLK (nx7631)
          ) ;
    nand02 ix4455 (.Y (nx4454), .A0 (nx5481), .A1 (nx7871)) ;
    nand03 ix5482 (.Y (nx5481), .A0 (nx5305), .A1 (nx7635), .A2 (nx4446)) ;
    nor02_2x ix4447 (.Y (nx4446), .A0 (nx4318), .A1 (nx4239)) ;
    nand02 ix4665 (.Y (nx4664), .A0 (nx5497), .A1 (nx7871)) ;
    nand03 ix5498 (.Y (nx5497), .A0 (nx5333), .A1 (nx7635), .A2 (nx4446)) ;
    latch i7_r15_lat_q_5 (.Q (DecompressedData1[109]), .D (nx7553), .CLK (nx7651
          )) ;
    latch i7_r15_lat_q_6 (.Q (DecompressedData1[110]), .D (nx7559), .CLK (nx7651
          )) ;
    latch i7_r15_lat_q_7 (.Q (DecompressedData1[111]), .D (nx7565), .CLK (nx7651
          )) ;
    nand02 ix4839 (.Y (nx4838), .A0 (nx5509), .A1 (nx7873)) ;
    nand03 ix5510 (.Y (nx5509), .A0 (nx5349), .A1 (nx7635), .A2 (nx4446)) ;
    nand02 ix5049 (.Y (nx5048), .A0 (nx5522), .A1 (nx7873)) ;
    nand03 ix5523 (.Y (nx5522), .A0 (nx7837), .A1 (nx7635), .A2 (nx4446)) ;
    latch i7_r13_lat_q_5 (.Q (DecompressedData1[125]), .D (nx7555), .CLK (nx7663
          )) ;
    latch i7_r13_lat_q_6 (.Q (DecompressedData1[126]), .D (nx7561), .CLK (nx7663
          )) ;
    latch i7_r13_lat_q_7 (.Q (DecompressedData1[127]), .D (nx7567), .CLK (nx7663
          )) ;
    nand02 ix5229 (.Y (nx5228), .A0 (nx5535), .A1 (nx7873)) ;
    nand03 ix5536 (.Y (nx5535), .A0 (nx5305), .A1 (nx7635), .A2 (nx5220)) ;
    nor02_2x ix5221 (.Y (nx5220), .A0 (nx4318), .A1 (i7_counterout2_2)) ;
    nand02 ix5447 (.Y (nx5446), .A0 (nx5549), .A1 (nx7873)) ;
    nand03 ix5550 (.Y (nx5549), .A0 (nx5333), .A1 (nx7635), .A2 (nx5220)) ;
    latch i7_r11_lat_q_5 (.Q (DecompressedData1[141]), .D (nx7555), .CLK (nx7675
          )) ;
    latch i7_r11_lat_q_6 (.Q (DecompressedData1[142]), .D (nx7561), .CLK (nx7675
          )) ;
    latch i7_r11_lat_q_7 (.Q (DecompressedData1[143]), .D (nx7567), .CLK (nx7675
          )) ;
    nand02 ix5621 (.Y (nx5620), .A0 (nx5562), .A1 (nx7873)) ;
    nand03 ix5563 (.Y (nx5562), .A0 (nx5349), .A1 (nx7637), .A2 (nx5220)) ;
    nand02 ix5831 (.Y (nx5830), .A0 (nx5576), .A1 (nx7873)) ;
    nand03 ix5577 (.Y (nx5576), .A0 (nx7837), .A1 (nx7637), .A2 (nx5220)) ;
    latch i7_r9_lat_q_5 (.Q (DecompressedData1[157]), .D (nx7555), .CLK (nx7687)
          ) ;
    latch i7_r9_lat_q_6 (.Q (DecompressedData1[158]), .D (nx7561), .CLK (nx7687)
          ) ;
    latch i7_r9_lat_q_7 (.Q (DecompressedData1[159]), .D (nx7567), .CLK (nx7687)
          ) ;
    nand02 ix6011 (.Y (nx6010), .A0 (nx5589), .A1 (nx7873)) ;
    nand03 ix5590 (.Y (nx5589), .A0 (nx5305), .A1 (nx7637), .A2 (nx6002)) ;
    nor02_2x ix6003 (.Y (nx6002), .A0 (i7_counterout2_3), .A1 (nx4239)) ;
    nand02 ix6221 (.Y (nx6220), .A0 (nx5603), .A1 (nx7875)) ;
    nand03 ix5604 (.Y (nx5603), .A0 (nx5333), .A1 (nx7637), .A2 (nx6002)) ;
    latch i7_r7_lat_q_5 (.Q (DecompressedData1[173]), .D (nx7555), .CLK (nx7699)
          ) ;
    latch i7_r7_lat_q_6 (.Q (DecompressedData1[174]), .D (nx7561), .CLK (nx7699)
          ) ;
    latch i7_r7_lat_q_7 (.Q (DecompressedData1[175]), .D (nx7567), .CLK (nx7699)
          ) ;
    nand02 ix6395 (.Y (nx6394), .A0 (nx5615), .A1 (nx7875)) ;
    nand03 ix5616 (.Y (nx5615), .A0 (nx5349), .A1 (nx7637), .A2 (nx6002)) ;
    nand02 ix6605 (.Y (nx6604), .A0 (nx5628), .A1 (nx7875)) ;
    nand03 ix5629 (.Y (nx5628), .A0 (nx4293), .A1 (nx7637), .A2 (nx6002)) ;
    latch i7_r5_lat_q_5 (.Q (DecompressedData1[189]), .D (nx7555), .CLK (nx7711)
          ) ;
    latch i7_r5_lat_q_6 (.Q (DecompressedData1[190]), .D (nx7561), .CLK (nx7711)
          ) ;
    latch i7_r5_lat_q_7 (.Q (DecompressedData1[191]), .D (nx7567), .CLK (nx7711)
          ) ;
    nand02 ix6787 (.Y (nx6786), .A0 (nx5643), .A1 (nx7875)) ;
    nand03 ix5644 (.Y (nx5643), .A0 (nx5305), .A1 (nx7639), .A2 (nx6778)) ;
    nor02_2x ix6779 (.Y (nx6778), .A0 (i7_counterout2_3), .A1 (i7_counterout2_2)
             ) ;
    nand02 ix6997 (.Y (nx6996), .A0 (nx5659), .A1 (nx7875)) ;
    nand03 ix5660 (.Y (nx5659), .A0 (nx5333), .A1 (nx7639), .A2 (nx6778)) ;
    latch i7_r3_lat_q_5 (.Q (DecompressedData1[205]), .D (nx7555), .CLK (nx7723)
          ) ;
    latch i7_r3_lat_q_6 (.Q (DecompressedData1[206]), .D (nx7561), .CLK (nx7723)
          ) ;
    latch i7_r3_lat_q_7 (.Q (DecompressedData1[207]), .D (nx7567), .CLK (nx7723)
          ) ;
    nand02 ix7171 (.Y (nx7170), .A0 (nx5671), .A1 (nx7875)) ;
    nand03 ix5672 (.Y (nx5671), .A0 (nx5349), .A1 (nx7639), .A2 (nx6778)) ;
    nand02 ix7381 (.Y (nx7380), .A0 (nx5684), .A1 (nx7875)) ;
    nand03 ix5685 (.Y (nx5684), .A0 (nx4293), .A1 (nx7639), .A2 (nx6778)) ;
    latch i7_r1_lat_q_5 (.Q (DecompressedData1[221]), .D (nx7555), .CLK (nx7735)
          ) ;
    latch i7_r1_lat_q_6 (.Q (DecompressedData1[222]), .D (nx7561), .CLK (nx7735)
          ) ;
    latch i7_r1_lat_q_7 (.Q (DecompressedData1[223]), .D (nx7567), .CLK (nx7735)
          ) ;
    mux21 ix2133 (.Y (DecompressedData[0]), .A0 (nx5695), .A1 (nx5697), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2159 (.Y (DecompressedData[1]), .A0 (nx5700), .A1 (nx5703), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2185 (.Y (DecompressedData[2]), .A0 (nx5707), .A1 (nx5709), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2211 (.Y (DecompressedData[3]), .A0 (nx5712), .A1 (nx5715), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2237 (.Y (DecompressedData[4]), .A0 (nx5719), .A1 (nx5721), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2263 (.Y (DecompressedData[5]), .A0 (nx5724), .A1 (nx5727), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2289 (.Y (DecompressedData[6]), .A0 (nx5731), .A1 (nx5733), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2315 (.Y (DecompressedData[7]), .A0 (nx5736), .A1 (nx5739), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2345 (.Y (DecompressedData[8]), .A0 (nx5743), .A1 (nx5745), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2369 (.Y (DecompressedData[9]), .A0 (nx5748), .A1 (nx5751), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2393 (.Y (DecompressedData[10]), .A0 (nx5755), .A1 (nx5757), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2417 (.Y (DecompressedData[11]), .A0 (nx5760), .A1 (nx5763), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2441 (.Y (DecompressedData[12]), .A0 (nx5767), .A1 (nx5769), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix2465 (.Y (DecompressedData[13]), .A0 (nx5772), .A1 (nx5775)) ;
    nand02 ix5773 (.Y (nx5772), .A0 (nx7743), .A1 (DecompressedData1[13])) ;
    nand02 ix5776 (.Y (nx5775), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[15])) ;
    nand02 ix2477 (.Y (DecompressedData[14]), .A0 (nx5779), .A1 (nx5775)) ;
    nand02 ix5780 (.Y (nx5779), .A0 (nx7743), .A1 (DecompressedData1[14])) ;
    nand02 ix2489 (.Y (DecompressedData[15]), .A0 (nx5782), .A1 (nx5775)) ;
    nand02 ix5783 (.Y (nx5782), .A0 (nx7743), .A1 (DecompressedData1[15])) ;
    mux21 ix2535 (.Y (DecompressedData[16]), .A0 (nx5785), .A1 (nx5787), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2559 (.Y (DecompressedData[17]), .A0 (nx5791), .A1 (nx5793), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2583 (.Y (DecompressedData[18]), .A0 (nx5796), .A1 (nx5799), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2607 (.Y (DecompressedData[19]), .A0 (nx5803), .A1 (nx5805), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2631 (.Y (DecompressedData[20]), .A0 (nx5808), .A1 (nx5811), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2655 (.Y (DecompressedData[21]), .A0 (nx5815), .A1 (nx5817), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2679 (.Y (DecompressedData[22]), .A0 (nx5820), .A1 (nx5823), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2703 (.Y (DecompressedData[23]), .A0 (nx5827), .A1 (nx5829), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2733 (.Y (DecompressedData[24]), .A0 (nx5833), .A1 (nx5835), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2757 (.Y (DecompressedData[25]), .A0 (nx5838), .A1 (nx5841), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2781 (.Y (DecompressedData[26]), .A0 (nx5845), .A1 (nx5847), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2805 (.Y (DecompressedData[27]), .A0 (nx5850), .A1 (nx5853), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2829 (.Y (DecompressedData[28]), .A0 (nx5857), .A1 (nx5859), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix2853 (.Y (DecompressedData[29]), .A0 (nx5862), .A1 (nx5865)) ;
    nand02 ix5863 (.Y (nx5862), .A0 (nx7743), .A1 (DecompressedData1[29])) ;
    nand02 ix5866 (.Y (nx5865), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[31])) ;
    nand02 ix2865 (.Y (DecompressedData[30]), .A0 (nx5869), .A1 (nx5865)) ;
    nand02 ix5870 (.Y (nx5869), .A0 (nx7743), .A1 (DecompressedData1[30])) ;
    nand02 ix2877 (.Y (DecompressedData[31]), .A0 (nx5872), .A1 (nx5865)) ;
    nand02 ix5873 (.Y (nx5872), .A0 (nx7743), .A1 (DecompressedData1[31])) ;
    mux21 ix2925 (.Y (DecompressedData[32]), .A0 (nx5875), .A1 (nx5877), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2949 (.Y (DecompressedData[33]), .A0 (nx5881), .A1 (nx5883), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2973 (.Y (DecompressedData[34]), .A0 (nx5886), .A1 (nx5889), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix2997 (.Y (DecompressedData[35]), .A0 (nx5893), .A1 (nx5895), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3021 (.Y (DecompressedData[36]), .A0 (nx5898), .A1 (nx5901), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3045 (.Y (DecompressedData[37]), .A0 (nx5905), .A1 (nx5907), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3069 (.Y (DecompressedData[38]), .A0 (nx5910), .A1 (nx5913), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3093 (.Y (DecompressedData[39]), .A0 (nx5917), .A1 (nx5919), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3123 (.Y (DecompressedData[40]), .A0 (nx5922), .A1 (nx5925), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3147 (.Y (DecompressedData[41]), .A0 (nx5929), .A1 (nx5931), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3171 (.Y (DecompressedData[42]), .A0 (nx5934), .A1 (nx5937), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3195 (.Y (DecompressedData[43]), .A0 (nx5941), .A1 (nx5943), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3219 (.Y (DecompressedData[44]), .A0 (nx5946), .A1 (nx5949), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix3243 (.Y (DecompressedData[45]), .A0 (nx5953), .A1 (nx5955)) ;
    nand02 ix5954 (.Y (nx5953), .A0 (nx7745), .A1 (DecompressedData1[45])) ;
    nand02 ix5956 (.Y (nx5955), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[47])) ;
    nand02 ix3255 (.Y (DecompressedData[46]), .A0 (nx5958), .A1 (nx5955)) ;
    nand02 ix5959 (.Y (nx5958), .A0 (nx7745), .A1 (DecompressedData1[46])) ;
    nand02 ix3267 (.Y (DecompressedData[47]), .A0 (nx5961), .A1 (nx5955)) ;
    nand02 ix5962 (.Y (nx5961), .A0 (nx7745), .A1 (DecompressedData1[47])) ;
    mux21 ix3313 (.Y (DecompressedData[48]), .A0 (nx5965), .A1 (nx5967), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3337 (.Y (DecompressedData[49]), .A0 (nx5970), .A1 (nx5973), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3361 (.Y (DecompressedData[50]), .A0 (nx5977), .A1 (nx5979), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3385 (.Y (DecompressedData[51]), .A0 (nx5982), .A1 (nx5985), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3409 (.Y (DecompressedData[52]), .A0 (nx5989), .A1 (nx5991), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3433 (.Y (DecompressedData[53]), .A0 (nx5994), .A1 (nx5997), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3457 (.Y (DecompressedData[54]), .A0 (nx6001), .A1 (nx6003), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3481 (.Y (DecompressedData[55]), .A0 (nx6007), .A1 (nx6009), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3511 (.Y (DecompressedData[56]), .A0 (nx6013), .A1 (nx6015), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3535 (.Y (DecompressedData[57]), .A0 (nx6018), .A1 (nx6021), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3559 (.Y (DecompressedData[58]), .A0 (nx6025), .A1 (nx6027), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3583 (.Y (DecompressedData[59]), .A0 (nx6031), .A1 (nx6033), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3607 (.Y (DecompressedData[60]), .A0 (nx6037), .A1 (nx6039), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix3631 (.Y (DecompressedData[61]), .A0 (nx6042), .A1 (nx6045)) ;
    nand02 ix6043 (.Y (nx6042), .A0 (nx7745), .A1 (DecompressedData1[61])) ;
    nand02 ix6046 (.Y (nx6045), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[63])) ;
    nand02 ix3643 (.Y (DecompressedData[62]), .A0 (nx6049), .A1 (nx6045)) ;
    nand02 ix6050 (.Y (nx6049), .A0 (nx7745), .A1 (DecompressedData1[62])) ;
    nand02 ix3655 (.Y (DecompressedData[63]), .A0 (nx6052), .A1 (nx6045)) ;
    nand02 ix6053 (.Y (nx6052), .A0 (nx7745), .A1 (DecompressedData1[63])) ;
    mux21 ix3713 (.Y (DecompressedData[64]), .A0 (nx6055), .A1 (nx6057), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3737 (.Y (DecompressedData[65]), .A0 (nx6061), .A1 (nx6063), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3761 (.Y (DecompressedData[66]), .A0 (nx6066), .A1 (nx6069), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3785 (.Y (DecompressedData[67]), .A0 (nx6073), .A1 (nx6075), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3809 (.Y (DecompressedData[68]), .A0 (nx6078), .A1 (nx6081), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3833 (.Y (DecompressedData[69]), .A0 (nx6085), .A1 (nx6087), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3857 (.Y (DecompressedData[70]), .A0 (nx6090), .A1 (nx6093), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3881 (.Y (DecompressedData[71]), .A0 (nx6097), .A1 (nx6099), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3911 (.Y (DecompressedData[72]), .A0 (nx6102), .A1 (nx6105), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3935 (.Y (DecompressedData[73]), .A0 (nx6109), .A1 (nx6111), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3959 (.Y (DecompressedData[74]), .A0 (nx6114), .A1 (nx6117), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix3983 (.Y (DecompressedData[75]), .A0 (nx6121), .A1 (nx6123), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4007 (.Y (DecompressedData[76]), .A0 (nx6126), .A1 (nx6129), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix4031 (.Y (DecompressedData[77]), .A0 (nx6133), .A1 (nx6135)) ;
    nand02 ix6134 (.Y (nx6133), .A0 (nx7745), .A1 (DecompressedData1[77])) ;
    nand02 ix6136 (.Y (nx6135), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[79])) ;
    nand02 ix4043 (.Y (DecompressedData[78]), .A0 (nx6138), .A1 (nx6135)) ;
    nand02 ix6139 (.Y (nx6138), .A0 (nx7747), .A1 (DecompressedData1[78])) ;
    nand02 ix4055 (.Y (DecompressedData[79]), .A0 (nx6141), .A1 (nx6135)) ;
    nand02 ix6142 (.Y (nx6141), .A0 (nx7747), .A1 (DecompressedData1[79])) ;
    mux21 ix4097 (.Y (DecompressedData[80]), .A0 (nx6145), .A1 (nx6147), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4121 (.Y (DecompressedData[81]), .A0 (nx6150), .A1 (nx6153), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4145 (.Y (DecompressedData[82]), .A0 (nx6157), .A1 (nx6159), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4169 (.Y (DecompressedData[83]), .A0 (nx6162), .A1 (nx6165), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4193 (.Y (DecompressedData[84]), .A0 (nx6169), .A1 (nx6171), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4217 (.Y (DecompressedData[85]), .A0 (nx6174), .A1 (nx6177), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4241 (.Y (DecompressedData[86]), .A0 (nx6181), .A1 (nx6183), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4265 (.Y (DecompressedData[87]), .A0 (nx6186), .A1 (nx6189), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4295 (.Y (DecompressedData[88]), .A0 (nx6193), .A1 (nx6195), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4319 (.Y (DecompressedData[89]), .A0 (nx6198), .A1 (nx6201), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4343 (.Y (DecompressedData[90]), .A0 (nx6205), .A1 (nx6207), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4367 (.Y (DecompressedData[91]), .A0 (nx6210), .A1 (nx6213), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4391 (.Y (DecompressedData[92]), .A0 (nx6217), .A1 (nx6219), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix4415 (.Y (DecompressedData[93]), .A0 (nx6223), .A1 (nx6225)) ;
    nand02 ix6224 (.Y (nx6223), .A0 (nx7747), .A1 (DecompressedData1[93])) ;
    nand02 ix6226 (.Y (nx6225), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[95])) ;
    nand02 ix4427 (.Y (DecompressedData[94]), .A0 (nx6228), .A1 (nx6225)) ;
    nand02 ix6229 (.Y (nx6228), .A0 (nx7747), .A1 (DecompressedData1[94])) ;
    nand02 ix4439 (.Y (DecompressedData[95]), .A0 (nx6231), .A1 (nx6225)) ;
    nand02 ix6232 (.Y (nx6231), .A0 (nx7747), .A1 (DecompressedData1[95])) ;
    mux21 ix4491 (.Y (DecompressedData[96]), .A0 (nx6235), .A1 (nx6237), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4515 (.Y (DecompressedData[97]), .A0 (nx6240), .A1 (nx6243), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4539 (.Y (DecompressedData[98]), .A0 (nx6247), .A1 (nx6249), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4563 (.Y (DecompressedData[99]), .A0 (nx6252), .A1 (nx6255), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4587 (.Y (DecompressedData[100]), .A0 (nx6259), .A1 (nx6261), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4611 (.Y (DecompressedData[101]), .A0 (nx6264), .A1 (nx6267), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4635 (.Y (DecompressedData[102]), .A0 (nx6271), .A1 (nx6273), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4659 (.Y (DecompressedData[103]), .A0 (nx6276), .A1 (nx6279), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4689 (.Y (DecompressedData[104]), .A0 (nx6283), .A1 (nx6285), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4713 (.Y (DecompressedData[105]), .A0 (nx6288), .A1 (nx6291), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4737 (.Y (DecompressedData[106]), .A0 (nx6295), .A1 (nx6297), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4761 (.Y (DecompressedData[107]), .A0 (nx6300), .A1 (nx6303), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4785 (.Y (DecompressedData[108]), .A0 (nx6307), .A1 (nx6309), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix4809 (.Y (DecompressedData[109]), .A0 (nx6312), .A1 (nx6315)) ;
    nand02 ix6313 (.Y (nx6312), .A0 (nx7747), .A1 (DecompressedData1[109])) ;
    nand02 ix6316 (.Y (nx6315), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[111])
           ) ;
    nand02 ix4821 (.Y (DecompressedData[110]), .A0 (nx6319), .A1 (nx6315)) ;
    nand02 ix6320 (.Y (nx6319), .A0 (nx7747), .A1 (DecompressedData1[110])) ;
    nand02 ix4833 (.Y (DecompressedData[111]), .A0 (nx6322), .A1 (nx6315)) ;
    nand02 ix6323 (.Y (nx6322), .A0 (nx7749), .A1 (DecompressedData1[111])) ;
    mux21 ix4875 (.Y (DecompressedData[112]), .A0 (nx6325), .A1 (nx6327), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4899 (.Y (DecompressedData[113]), .A0 (nx6331), .A1 (nx6333), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4923 (.Y (DecompressedData[114]), .A0 (nx6336), .A1 (nx6339), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4947 (.Y (DecompressedData[115]), .A0 (nx6343), .A1 (nx6345), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4971 (.Y (DecompressedData[116]), .A0 (nx6348), .A1 (nx6350), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix4995 (.Y (DecompressedData[117]), .A0 (nx6353), .A1 (nx6355), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5019 (.Y (DecompressedData[118]), .A0 (nx6358), .A1 (nx6360), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5043 (.Y (DecompressedData[119]), .A0 (nx6363), .A1 (nx6365), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5073 (.Y (DecompressedData[120]), .A0 (nx6368), .A1 (nx6370), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5097 (.Y (DecompressedData[121]), .A0 (nx6373), .A1 (nx6375), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5121 (.Y (DecompressedData[122]), .A0 (nx6379), .A1 (nx6381), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5145 (.Y (DecompressedData[123]), .A0 (nx6384), .A1 (nx6387), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5169 (.Y (DecompressedData[124]), .A0 (nx6391), .A1 (nx6393), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix5193 (.Y (DecompressedData[125]), .A0 (nx6397), .A1 (nx6399)) ;
    nand02 ix6398 (.Y (nx6397), .A0 (nx7749), .A1 (DecompressedData1[125])) ;
    nand02 ix6400 (.Y (nx6399), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[127])
           ) ;
    nand02 ix5205 (.Y (DecompressedData[126]), .A0 (nx6402), .A1 (nx6399)) ;
    nand02 ix6403 (.Y (nx6402), .A0 (nx7749), .A1 (DecompressedData1[126])) ;
    nand02 ix5217 (.Y (DecompressedData[127]), .A0 (nx6405), .A1 (nx6399)) ;
    nand02 ix6406 (.Y (nx6405), .A0 (nx7749), .A1 (DecompressedData1[127])) ;
    mux21 ix5273 (.Y (DecompressedData[128]), .A0 (nx6409), .A1 (nx6411), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5297 (.Y (DecompressedData[129]), .A0 (nx6415), .A1 (nx6417), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5321 (.Y (DecompressedData[130]), .A0 (nx6421), .A1 (nx6423), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5345 (.Y (DecompressedData[131]), .A0 (nx6426), .A1 (nx6429), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5369 (.Y (DecompressedData[132]), .A0 (nx6433), .A1 (nx6435), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5393 (.Y (DecompressedData[133]), .A0 (nx6438), .A1 (nx6441), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5417 (.Y (DecompressedData[134]), .A0 (nx6445), .A1 (nx6447), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5441 (.Y (DecompressedData[135]), .A0 (nx6450), .A1 (nx6453), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5471 (.Y (DecompressedData[136]), .A0 (nx6457), .A1 (nx6459), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5495 (.Y (DecompressedData[137]), .A0 (nx6462), .A1 (nx6465), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5519 (.Y (DecompressedData[138]), .A0 (nx6469), .A1 (nx6471), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5543 (.Y (DecompressedData[139]), .A0 (nx6474), .A1 (nx6477), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5567 (.Y (DecompressedData[140]), .A0 (nx6481), .A1 (nx6483), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix5591 (.Y (DecompressedData[141]), .A0 (nx6486), .A1 (nx6489)) ;
    nand02 ix6487 (.Y (nx6486), .A0 (nx7749), .A1 (DecompressedData1[141])) ;
    nand02 ix6490 (.Y (nx6489), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[143])
           ) ;
    nand02 ix5603 (.Y (DecompressedData[142]), .A0 (nx6493), .A1 (nx6489)) ;
    nand02 ix6494 (.Y (nx6493), .A0 (nx7749), .A1 (DecompressedData1[142])) ;
    nand02 ix5615 (.Y (DecompressedData[143]), .A0 (nx6496), .A1 (nx6489)) ;
    nand02 ix6497 (.Y (nx6496), .A0 (nx7749), .A1 (DecompressedData1[143])) ;
    mux21 ix5657 (.Y (DecompressedData[144]), .A0 (nx6499), .A1 (nx6501), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5681 (.Y (DecompressedData[145]), .A0 (nx6505), .A1 (nx6507), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5705 (.Y (DecompressedData[146]), .A0 (nx6510), .A1 (nx6513), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5729 (.Y (DecompressedData[147]), .A0 (nx6517), .A1 (nx6519), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5753 (.Y (DecompressedData[148]), .A0 (nx6522), .A1 (nx6525), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5777 (.Y (DecompressedData[149]), .A0 (nx6529), .A1 (nx6531), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5801 (.Y (DecompressedData[150]), .A0 (nx6534), .A1 (nx6537), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5825 (.Y (DecompressedData[151]), .A0 (nx6541), .A1 (nx6543), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5855 (.Y (DecompressedData[152]), .A0 (nx6546), .A1 (nx6549), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5879 (.Y (DecompressedData[153]), .A0 (nx6553), .A1 (nx6555), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5903 (.Y (DecompressedData[154]), .A0 (nx6558), .A1 (nx6561), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5927 (.Y (DecompressedData[155]), .A0 (nx6565), .A1 (nx6567), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix5951 (.Y (DecompressedData[156]), .A0 (nx6570), .A1 (nx6573), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix5975 (.Y (DecompressedData[157]), .A0 (nx6577), .A1 (nx6579)) ;
    nand02 ix6578 (.Y (nx6577), .A0 (nx7751), .A1 (DecompressedData1[157])) ;
    nand02 ix6580 (.Y (nx6579), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[159])
           ) ;
    nand02 ix5987 (.Y (DecompressedData[158]), .A0 (nx6582), .A1 (nx6579)) ;
    nand02 ix6583 (.Y (nx6582), .A0 (nx7751), .A1 (DecompressedData1[158])) ;
    nand02 ix5999 (.Y (DecompressedData[159]), .A0 (nx6585), .A1 (nx6579)) ;
    nand02 ix6586 (.Y (nx6585), .A0 (nx7751), .A1 (DecompressedData1[159])) ;
    mux21 ix6047 (.Y (DecompressedData[160]), .A0 (nx6589), .A1 (nx6591), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6071 (.Y (DecompressedData[161]), .A0 (nx6594), .A1 (nx6597), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6095 (.Y (DecompressedData[162]), .A0 (nx6601), .A1 (nx6603), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6119 (.Y (DecompressedData[163]), .A0 (nx6607), .A1 (nx6609), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6143 (.Y (DecompressedData[164]), .A0 (nx6612), .A1 (nx6615), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6167 (.Y (DecompressedData[165]), .A0 (nx6619), .A1 (nx6621), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6191 (.Y (DecompressedData[166]), .A0 (nx6624), .A1 (nx6627), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6215 (.Y (DecompressedData[167]), .A0 (nx6631), .A1 (nx6633), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6245 (.Y (DecompressedData[168]), .A0 (nx6636), .A1 (nx6639), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6269 (.Y (DecompressedData[169]), .A0 (nx6643), .A1 (nx6645), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6293 (.Y (DecompressedData[170]), .A0 (nx6648), .A1 (nx6651), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6317 (.Y (DecompressedData[171]), .A0 (nx6655), .A1 (nx6657), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6341 (.Y (DecompressedData[172]), .A0 (nx6660), .A1 (nx6663), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix6365 (.Y (DecompressedData[173]), .A0 (nx6667), .A1 (nx6669)) ;
    nand02 ix6668 (.Y (nx6667), .A0 (nx7751), .A1 (DecompressedData1[173])) ;
    nand02 ix6670 (.Y (nx6669), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[175])
           ) ;
    nand02 ix6377 (.Y (DecompressedData[174]), .A0 (nx6672), .A1 (nx6669)) ;
    nand02 ix6673 (.Y (nx6672), .A0 (nx7751), .A1 (DecompressedData1[174])) ;
    nand02 ix6389 (.Y (DecompressedData[175]), .A0 (nx6675), .A1 (nx6669)) ;
    nand02 ix6676 (.Y (nx6675), .A0 (nx7751), .A1 (DecompressedData1[175])) ;
    mux21 ix6431 (.Y (DecompressedData[176]), .A0 (nx6679), .A1 (nx6681), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6455 (.Y (DecompressedData[177]), .A0 (nx6684), .A1 (nx6687), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6479 (.Y (DecompressedData[178]), .A0 (nx6691), .A1 (nx6693), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6503 (.Y (DecompressedData[179]), .A0 (nx6696), .A1 (nx6699), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6527 (.Y (DecompressedData[180]), .A0 (nx6703), .A1 (nx6705), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6551 (.Y (DecompressedData[181]), .A0 (nx6708), .A1 (nx6711), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6575 (.Y (DecompressedData[182]), .A0 (nx6715), .A1 (nx6717), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6599 (.Y (DecompressedData[183]), .A0 (nx6720), .A1 (nx6723), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6629 (.Y (DecompressedData[184]), .A0 (nx6727), .A1 (nx6729), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6653 (.Y (DecompressedData[185]), .A0 (nx6732), .A1 (nx6734), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6677 (.Y (DecompressedData[186]), .A0 (nx6737), .A1 (nx6739), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6701 (.Y (DecompressedData[187]), .A0 (nx6742), .A1 (nx6744), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6725 (.Y (DecompressedData[188]), .A0 (nx6747), .A1 (nx6749), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix6749 (.Y (DecompressedData[189]), .A0 (nx6752), .A1 (nx6754)) ;
    nand02 ix6753 (.Y (nx6752), .A0 (nx7751), .A1 (DecompressedData1[189])) ;
    nand02 ix6755 (.Y (nx6754), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[191])
           ) ;
    nand02 ix6761 (.Y (DecompressedData[190]), .A0 (nx6757), .A1 (nx6754)) ;
    nand02 ix6758 (.Y (nx6757), .A0 (nx7753), .A1 (DecompressedData1[190])) ;
    nand02 ix6773 (.Y (DecompressedData[191]), .A0 (nx6761), .A1 (nx6754)) ;
    nand02 ix6762 (.Y (nx6761), .A0 (nx7753), .A1 (DecompressedData1[191])) ;
    mux21 ix6823 (.Y (DecompressedData[192]), .A0 (nx6764), .A1 (nx6766), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6847 (.Y (DecompressedData[193]), .A0 (nx6769), .A1 (nx6771), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6871 (.Y (DecompressedData[194]), .A0 (nx6775), .A1 (nx6777), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6895 (.Y (DecompressedData[195]), .A0 (nx6781), .A1 (nx6783), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6919 (.Y (DecompressedData[196]), .A0 (nx6787), .A1 (nx6789), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6943 (.Y (DecompressedData[197]), .A0 (nx6792), .A1 (nx6794), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6967 (.Y (DecompressedData[198]), .A0 (nx6797), .A1 (nx6799), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix6991 (.Y (DecompressedData[199]), .A0 (nx6803), .A1 (nx6805), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7021 (.Y (DecompressedData[200]), .A0 (nx6809), .A1 (nx6811), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7045 (.Y (DecompressedData[201]), .A0 (nx6815), .A1 (nx6817), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7069 (.Y (DecompressedData[202]), .A0 (nx6821), .A1 (nx6823), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7093 (.Y (DecompressedData[203]), .A0 (nx6826), .A1 (nx6828), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7117 (.Y (DecompressedData[204]), .A0 (nx6831), .A1 (nx6833), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix7141 (.Y (DecompressedData[205]), .A0 (nx6837), .A1 (nx6839)) ;
    nand02 ix6838 (.Y (nx6837), .A0 (nx7753), .A1 (DecompressedData1[205])) ;
    nand02 ix6840 (.Y (nx6839), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[207])
           ) ;
    nand02 ix7153 (.Y (DecompressedData[206]), .A0 (nx6842), .A1 (nx6839)) ;
    nand02 ix6843 (.Y (nx6842), .A0 (nx7753), .A1 (DecompressedData1[206])) ;
    nand02 ix7165 (.Y (DecompressedData[207]), .A0 (nx6845), .A1 (nx6839)) ;
    nand02 ix6846 (.Y (nx6845), .A0 (nx7753), .A1 (DecompressedData1[207])) ;
    mux21 ix7207 (.Y (DecompressedData[208]), .A0 (nx6849), .A1 (nx6851), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7231 (.Y (DecompressedData[209]), .A0 (nx6854), .A1 (nx6857), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7255 (.Y (DecompressedData[210]), .A0 (nx6861), .A1 (nx6863), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7279 (.Y (DecompressedData[211]), .A0 (nx6866), .A1 (nx6869), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7303 (.Y (DecompressedData[212]), .A0 (nx6873), .A1 (nx6875), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7327 (.Y (DecompressedData[213]), .A0 (nx6878), .A1 (nx6881), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7351 (.Y (DecompressedData[214]), .A0 (nx6885), .A1 (nx6887), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7375 (.Y (DecompressedData[215]), .A0 (nx6890), .A1 (nx6893), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7405 (.Y (DecompressedData[216]), .A0 (nx6897), .A1 (nx6899), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7429 (.Y (DecompressedData[217]), .A0 (nx6902), .A1 (nx6905), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7453 (.Y (DecompressedData[218]), .A0 (nx6909), .A1 (nx6911), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7477 (.Y (DecompressedData[219]), .A0 (nx6914), .A1 (nx6917), .S0 (
          CNNIMGLOAD)) ;
    mux21 ix7501 (.Y (DecompressedData[220]), .A0 (nx6921), .A1 (nx6923), .S0 (
          CNNIMGLOAD)) ;
    nand02 ix7525 (.Y (DecompressedData[221]), .A0 (nx6926), .A1 (nx6929)) ;
    nand02 ix6927 (.Y (nx6926), .A0 (nx7753), .A1 (DecompressedData1[221])) ;
    nand02 ix6930 (.Y (nx6929), .A0 (CNNIMGLOAD), .A1 (DecompressedData2[223])
           ) ;
    nand02 ix7537 (.Y (DecompressedData[222]), .A0 (nx6933), .A1 (nx6929)) ;
    nand02 ix6934 (.Y (nx6933), .A0 (nx7753), .A1 (DecompressedData1[222])) ;
    nand02 ix7549 (.Y (DecompressedData[223]), .A0 (nx6936), .A1 (nx6929)) ;
    nand02 ix6937 (.Y (nx6936), .A0 (nx7755), .A1 (DecompressedData1[223])) ;
    nor02_2x ix1201 (.Y (DecompressedData[224]), .A0 (nx7755), .A1 (nx6939)) ;
    nor02_2x ix1215 (.Y (DecompressedData[225]), .A0 (nx7755), .A1 (nx6943)) ;
    nor02_2x ix1229 (.Y (DecompressedData[226]), .A0 (nx7755), .A1 (nx6946)) ;
    nor02_2x ix1243 (.Y (DecompressedData[227]), .A0 (nx7755), .A1 (nx6949)) ;
    nor02_2x ix1257 (.Y (DecompressedData[228]), .A0 (nx7755), .A1 (nx6953)) ;
    nor02_2x ix1271 (.Y (DecompressedData[229]), .A0 (nx7755), .A1 (nx6957)) ;
    nor02_2x ix1285 (.Y (DecompressedData[230]), .A0 (nx7757), .A1 (nx6960)) ;
    nor02_2x ix1299 (.Y (DecompressedData[231]), .A0 (nx7757), .A1 (nx6963)) ;
    nor02_2x ix1313 (.Y (DecompressedData[232]), .A0 (nx7757), .A1 (nx6967)) ;
    nor02_2x ix1327 (.Y (DecompressedData[233]), .A0 (nx7757), .A1 (nx6970)) ;
    nor02_2x ix1341 (.Y (DecompressedData[234]), .A0 (nx7757), .A1 (nx6973)) ;
    nor02_2x ix1355 (.Y (DecompressedData[235]), .A0 (nx7757), .A1 (nx6977)) ;
    nor02_2x ix1369 (.Y (DecompressedData[236]), .A0 (nx7757), .A1 (nx6981)) ;
    nor02_2x ix1383 (.Y (DecompressedData[239]), .A0 (nx7759), .A1 (nx6984)) ;
    nor02_2x ix1407 (.Y (DecompressedData[240]), .A0 (nx7759), .A1 (nx6987)) ;
    nor02_2x ix1419 (.Y (DecompressedData[241]), .A0 (nx7759), .A1 (nx6991)) ;
    nor02_2x ix1431 (.Y (DecompressedData[242]), .A0 (nx7759), .A1 (nx6995)) ;
    nor02_2x ix1443 (.Y (DecompressedData[243]), .A0 (nx7759), .A1 (nx6999)) ;
    nor02_2x ix1455 (.Y (DecompressedData[244]), .A0 (nx7759), .A1 (nx7002)) ;
    nor02_2x ix1467 (.Y (DecompressedData[245]), .A0 (nx7759), .A1 (nx7005)) ;
    nor02_2x ix1479 (.Y (DecompressedData[246]), .A0 (nx7761), .A1 (nx7009)) ;
    nor02_2x ix1491 (.Y (DecompressedData[247]), .A0 (nx7761), .A1 (nx7013)) ;
    nor02_2x ix1503 (.Y (DecompressedData[248]), .A0 (nx7761), .A1 (nx7016)) ;
    nor02_2x ix1515 (.Y (DecompressedData[249]), .A0 (nx7761), .A1 (nx7019)) ;
    nor02_2x ix1527 (.Y (DecompressedData[250]), .A0 (nx7761), .A1 (nx7023)) ;
    nor02_2x ix1539 (.Y (DecompressedData[251]), .A0 (nx7761), .A1 (nx7026)) ;
    nor02_2x ix1551 (.Y (DecompressedData[252]), .A0 (nx7761), .A1 (nx7029)) ;
    nor02_2x ix1563 (.Y (DecompressedData[255]), .A0 (nx7763), .A1 (nx7033)) ;
    inv01 ix7038 (.Y (nx7037), .A (OuterAddress[0])) ;
    dff i5_aa_reg_Q (.Q (i5_FAEN), .QB (\$dummy [10]), .D (nx1616), .CLK (CLK)
        ) ;
    nor02ii ix1617 (.Y (nx1616), .A0 (nx7045), .A1 (nx1614)) ;
    nor02_2x ix7046 (.Y (nx7045), .A0 (nx1606), .A1 (nx1604)) ;
    nor02_2x ix1607 (.Y (nx1606), .A0 (nx7957), .A1 (nx7048)) ;
    aoi21 ix7049 (.Y (nx7048), .A0 (OuterWrite), .A1 (ProcessEnable), .B0 (
          DecompressionDone)) ;
    nand02 ix1595 (.Y (DecompressionDone), .A0 (nx7051), .A1 (nx7057)) ;
    dffs_ni i7_reg_readtoRam (.Q (DecompressionDone1), .QB (nx7051), .D (nx3503)
            , .CLK (CLK), .S (NOT_nx814)) ;
    nor02_2x ix3504 (.Y (nx3503), .A0 (nx7051), .A1 (nx814)) ;
    dffs_ni i8_reg_ramWrite (.Q (DecompressionDone2), .QB (nx7057), .D (nx3493)
            , .CLK (CLK), .S (nx558)) ;
    nor02_2x ix3494 (.Y (nx3493), .A0 (nx7057), .A1 (nx546)) ;
    nand02 ix559 (.Y (nx558), .A0 (nx546), .A1 (nx4011)) ;
    nor03_2x ix1605 (.Y (nx1604), .A0 (nx3563), .A1 (nx7063), .A2 (nx1598)) ;
    inv01 ix7064 (.Y (nx7063), .A (INCEnable)) ;
    nand03 ix1599 (.Y (nx1598), .A0 (nx7067), .A1 (nx7051), .A2 (nx7057)) ;
    nand02 ix7068 (.Y (nx7067), .A0 (OuterWrite), .A1 (ProcessEnable)) ;
    nor02_2x ix1615 (.Y (nx1614), .A0 (Rst), .A1 (nx7515)) ;
    dffr i5_MR_reg_dataout_0 (.Q (i5_MARo_0), .QB (nx7039), .D (nx1634), .CLK (
         CLK), .R (Rst)) ;
    inv01 ix7080 (.Y (nx7079), .A (OuterAddress[1])) ;
    dffr i5_MR_reg_dataout_1 (.Q (i5_MARo_1), .QB (nx7081), .D (nx1660), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix1661 (.Y (nx1660), .A0 (nx7877), .A1 (nx7085), .B0 (nx7088)) ;
    xnor2 ix7086 (.Y (nx7085), .A0 (nx1626), .A1 (Address[1])) ;
    nand02 ix1627 (.Y (nx1626), .A0 (nx7072), .A1 (nx7515)) ;
    oai21 ix7089 (.Y (nx7088), .A0 (nx1670), .A1 (nx1668), .B0 (nx7877)) ;
    nor02_2x ix1671 (.Y (nx1670), .A0 (nx7079), .A1 (nx7889)) ;
    nor02_2x ix1669 (.Y (nx1668), .A0 (nx7081), .A1 (nx7521)) ;
    nor02_2x ix1643 (.Y (nx1642), .A0 (nx7095), .A1 (nx7907)) ;
    inv01 ix7096 (.Y (nx7095), .A (ActivateOuterAddress)) ;
    inv01 ix7099 (.Y (nx7098), .A (OuterAddress[2])) ;
    dffr i5_MR_reg_dataout_2 (.Q (i5_MARo_2), .QB (nx7100), .D (nx1688), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix1689 (.Y (nx1688), .A0 (nx7877), .A1 (nx7103), .B0 (nx7109)) ;
    xnor2 ix7104 (.Y (nx7103), .A0 (nx1682), .A1 (Address[2])) ;
    oai21 ix1683 (.Y (nx1682), .A0 (nx7072), .A1 (nx7107), .B0 (nx7515)) ;
    oai21 ix7110 (.Y (nx7109), .A0 (nx1698), .A1 (nx1696), .B0 (nx7877)) ;
    nor02_2x ix1699 (.Y (nx1698), .A0 (nx7098), .A1 (nx7889)) ;
    nor02_2x ix1697 (.Y (nx1696), .A0 (nx7100), .A1 (nx7521)) ;
    inv01 ix7116 (.Y (nx7115), .A (OuterAddress[3])) ;
    oai21 ix1717 (.Y (nx1716), .A0 (nx7877), .A1 (nx7121), .B0 (nx7132)) ;
    xnor2 ix7122 (.Y (nx7121), .A0 (nx7123), .A1 (nx7129)) ;
    nand02 ix7124 (.Y (nx7123), .A0 (nx1682), .A1 (nx1708)) ;
    nand02 ix1709 (.Y (nx1708), .A0 (nx7126), .A1 (nx7515)) ;
    dffr i5_MR_reg_dataout_3 (.Q (i5_MARo_3), .QB (nx7117), .D (nx1716), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7133 (.Y (nx7132), .A0 (nx1726), .A1 (nx1724), .B0 (nx7877)) ;
    nor02_2x ix1727 (.Y (nx1726), .A0 (nx7115), .A1 (nx7891)) ;
    nor02_2x ix1725 (.Y (nx1724), .A0 (nx7117), .A1 (nx7521)) ;
    inv01 ix7138 (.Y (nx7137), .A (OuterAddress[4])) ;
    oai21 ix1745 (.Y (nx1744), .A0 (nx7877), .A1 (nx7143), .B0 (nx7151)) ;
    xnor2 ix7144 (.Y (nx7143), .A0 (nx7145), .A1 (nx7148)) ;
    nand03 ix7146 (.Y (nx7145), .A0 (nx1682), .A1 (nx1708), .A2 (nx1736)) ;
    nand02 ix1737 (.Y (nx1736), .A0 (nx7129), .A1 (nx7515)) ;
    dffr i5_MR_reg_dataout_4 (.Q (i5_MARo_4), .QB (nx7139), .D (nx1744), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7152 (.Y (nx7151), .A0 (nx1754), .A1 (nx1752), .B0 (nx7879)) ;
    nor02_2x ix1755 (.Y (nx1754), .A0 (nx7137), .A1 (nx7891)) ;
    nor02_2x ix1753 (.Y (nx1752), .A0 (nx7139), .A1 (nx7521)) ;
    inv01 ix7158 (.Y (nx7157), .A (OuterAddress[5])) ;
    oai21 ix1773 (.Y (nx1772), .A0 (nx7879), .A1 (nx7163), .B0 (nx7173)) ;
    xnor2 ix7164 (.Y (nx7163), .A0 (nx7165), .A1 (nx7169)) ;
    nand04 ix7166 (.Y (nx7165), .A0 (nx1682), .A1 (nx1708), .A2 (nx1736), .A3 (
           nx1764)) ;
    nand02 ix1765 (.Y (nx1764), .A0 (nx7148), .A1 (nx7515)) ;
    dffr i5_MR_reg_dataout_5 (.Q (i5_MARo_5), .QB (nx7159), .D (nx1772), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7174 (.Y (nx7173), .A0 (nx1782), .A1 (nx1780), .B0 (nx7879)) ;
    nor02_2x ix1783 (.Y (nx1782), .A0 (nx7157), .A1 (nx7893)) ;
    nor02_2x ix1781 (.Y (nx1780), .A0 (nx7159), .A1 (nx7521)) ;
    inv01 ix7179 (.Y (nx7178), .A (OuterAddress[6])) ;
    dffr i5_MR_reg_dataout_6 (.Q (i5_MARo_6), .QB (nx7181), .D (nx1800), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix1801 (.Y (nx1800), .A0 (nx7879), .A1 (nx7185), .B0 (nx7189)) ;
    xnor2 ix7186 (.Y (nx7185), .A0 (nx7525), .A1 (Address[6])) ;
    aoi21 ix1795 (.Y (nx1794), .A0 (nx7169), .A1 (nx7517), .B0 (nx7165)) ;
    oai21 ix7190 (.Y (nx7189), .A0 (nx1810), .A1 (nx1808), .B0 (nx7879)) ;
    nor02_2x ix1811 (.Y (nx1810), .A0 (nx7178), .A1 (nx7893)) ;
    nor02_2x ix1809 (.Y (nx1808), .A0 (nx7181), .A1 (nx7521)) ;
    inv01 ix7198 (.Y (nx7197), .A (OuterAddress[7])) ;
    oai21 ix1829 (.Y (nx1828), .A0 (nx7879), .A1 (nx7202), .B0 (nx7214)) ;
    xnor2 ix7203 (.Y (nx7202), .A0 (nx7205), .A1 (nx7211)) ;
    nand02 ix7206 (.Y (nx7205), .A0 (nx7525), .A1 (nx1820)) ;
    nand02 ix1821 (.Y (nx1820), .A0 (nx7209), .A1 (nx7517)) ;
    dffr i5_MR_reg_dataout_7 (.Q (i5_MARo_7), .QB (nx7199), .D (nx1828), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7215 (.Y (nx7214), .A0 (nx1838), .A1 (nx1836), .B0 (nx7879)) ;
    nor02_2x ix1839 (.Y (nx1838), .A0 (nx7197), .A1 (nx7895)) ;
    nor02_2x ix1837 (.Y (nx1836), .A0 (nx7199), .A1 (nx7523)) ;
    inv01 ix7222 (.Y (nx7221), .A (OuterAddress[8])) ;
    oai21 ix1857 (.Y (nx1856), .A0 (nx7881), .A1 (nx7226), .B0 (nx7236)) ;
    xnor2 ix7227 (.Y (nx7226), .A0 (nx7229), .A1 (nx7233)) ;
    nand03 ix7230 (.Y (nx7229), .A0 (nx7525), .A1 (nx1820), .A2 (nx1848)) ;
    nand02 ix1849 (.Y (nx1848), .A0 (nx7211), .A1 (nx7517)) ;
    dffr i5_MR_reg_dataout_8 (.Q (i5_MARo_8), .QB (nx7223), .D (nx1856), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7237 (.Y (nx7236), .A0 (nx1866), .A1 (nx1864), .B0 (nx7881)) ;
    nor02_2x ix1867 (.Y (nx1866), .A0 (nx7221), .A1 (nx7895)) ;
    nor02_2x ix1865 (.Y (nx1864), .A0 (nx7223), .A1 (nx7523)) ;
    inv01 ix7242 (.Y (nx7241), .A (OuterAddress[9])) ;
    oai21 ix1885 (.Y (nx1884), .A0 (nx7881), .A1 (nx7247), .B0 (nx7257)) ;
    xnor2 ix7248 (.Y (nx7247), .A0 (nx7249), .A1 (nx7253)) ;
    nand04 ix7250 (.Y (nx7249), .A0 (nx7525), .A1 (nx1820), .A2 (nx1848), .A3 (
           nx1876)) ;
    nand02 ix1877 (.Y (nx1876), .A0 (nx7233), .A1 (nx7517)) ;
    dffr i5_MR_reg_dataout_9 (.Q (i5_MARo_9), .QB (nx7243), .D (nx1884), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7258 (.Y (nx7257), .A0 (nx1894), .A1 (nx1892), .B0 (nx7881)) ;
    nor02_2x ix1895 (.Y (nx1894), .A0 (nx7241), .A1 (nx7895)) ;
    nor02_2x ix1893 (.Y (nx1892), .A0 (nx7243), .A1 (nx7523)) ;
    inv01 ix7263 (.Y (nx7262), .A (OuterAddress[10])) ;
    dffr i5_MR_reg_dataout_10 (.Q (i5_MARo_10), .QB (nx7265), .D (nx1912), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix1913 (.Y (nx1912), .A0 (nx7881), .A1 (nx7269), .B0 (nx7272)) ;
    xnor2 ix7270 (.Y (nx7269), .A0 (nx7527), .A1 (Address[10])) ;
    aoi21 ix1907 (.Y (nx1906), .A0 (nx7253), .A1 (nx7517), .B0 (nx7249)) ;
    oai21 ix7273 (.Y (nx7272), .A0 (nx1922), .A1 (nx1920), .B0 (nx7881)) ;
    nor02_2x ix1923 (.Y (nx1922), .A0 (nx7262), .A1 (nx7897)) ;
    nor02_2x ix1921 (.Y (nx1920), .A0 (nx7265), .A1 (nx7523)) ;
    inv01 ix7278 (.Y (nx7277), .A (OuterAddress[11])) ;
    oai21 ix1941 (.Y (nx1940), .A0 (nx7881), .A1 (nx7282), .B0 (nx7293)) ;
    xnor2 ix7283 (.Y (nx7282), .A0 (nx7284), .A1 (nx7289)) ;
    nand02 ix7285 (.Y (nx7284), .A0 (nx7527), .A1 (nx1932)) ;
    nand02 ix1933 (.Y (nx1932), .A0 (nx7287), .A1 (nx7517)) ;
    dffr i5_MR_reg_dataout_11 (.Q (i5_MARo_11), .QB (nx7279), .D (nx1940), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7294 (.Y (nx7293), .A0 (nx1950), .A1 (nx1948), .B0 (nx7883)) ;
    nor02_2x ix1951 (.Y (nx1950), .A0 (nx7277), .A1 (nx7897)) ;
    nor02_2x ix1949 (.Y (nx1948), .A0 (nx7279), .A1 (nx7523)) ;
    inv01 ix7299 (.Y (nx7298), .A (OuterAddress[12])) ;
    oai21 ix1969 (.Y (nx1968), .A0 (nx7883), .A1 (nx7305), .B0 (nx7313)) ;
    xnor2 ix7306 (.Y (nx7305), .A0 (nx7307), .A1 (nx7310)) ;
    nand03 ix7308 (.Y (nx7307), .A0 (nx7527), .A1 (nx1932), .A2 (nx1960)) ;
    nand02 ix1961 (.Y (nx1960), .A0 (nx7289), .A1 (nx7517)) ;
    dffr i5_MR_reg_dataout_12 (.Q (i5_MARo_12), .QB (nx7301), .D (nx1968), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7314 (.Y (nx7313), .A0 (nx1978), .A1 (nx1976), .B0 (nx7883)) ;
    nor02_2x ix1979 (.Y (nx1978), .A0 (nx7298), .A1 (nx7899)) ;
    nor02_2x ix1977 (.Y (nx1976), .A0 (nx7301), .A1 (nx7523)) ;
    inv01 ix7320 (.Y (nx7319), .A (OuterAddress[13])) ;
    oai21 ix1997 (.Y (nx1996), .A0 (nx7883), .A1 (nx7325), .B0 (nx7333)) ;
    xnor2 ix7326 (.Y (nx7325), .A0 (nx7327), .A1 (nx7330)) ;
    nand04 ix7328 (.Y (nx7327), .A0 (nx7527), .A1 (nx1932), .A2 (nx1960), .A3 (
           nx1988)) ;
    nand02 ix1989 (.Y (nx1988), .A0 (nx7310), .A1 (nx7519)) ;
    dffr i5_MR_reg_dataout_13 (.Q (i5_MARo_13), .QB (nx7321), .D (nx1996), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7334 (.Y (nx7333), .A0 (nx2006), .A1 (nx2004), .B0 (nx7883)) ;
    nor02_2x ix2007 (.Y (nx2006), .A0 (nx7319), .A1 (nx7899)) ;
    nor02_2x ix2005 (.Y (nx2004), .A0 (nx7321), .A1 (nx1642)) ;
    inv01 ix7340 (.Y (nx7339), .A (OuterAddress[14])) ;
    dffr i5_MR_reg_dataout_14 (.Q (i5_MARo_14), .QB (nx7341), .D (nx2024), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix2025 (.Y (nx2024), .A0 (nx7883), .A1 (nx7344), .B0 (nx7347)) ;
    xnor2 ix7345 (.Y (nx7344), .A0 (nx2018), .A1 (Address[14])) ;
    aoi21 ix2019 (.Y (nx2018), .A0 (nx7330), .A1 (nx7519), .B0 (nx7327)) ;
    oai21 ix7348 (.Y (nx7347), .A0 (nx2034), .A1 (nx2032), .B0 (nx7883)) ;
    nor02_2x ix2035 (.Y (nx2034), .A0 (nx7339), .A1 (nx7899)) ;
    nor02_2x ix2033 (.Y (nx2032), .A0 (nx7341), .A1 (nx1642)) ;
    inv01 ix7355 (.Y (nx7354), .A (OuterAddress[15])) ;
    oai21 ix2053 (.Y (nx2052), .A0 (nx7885), .A1 (nx7359), .B0 (nx7370)) ;
    xnor2 ix7360 (.Y (nx7359), .A0 (nx7361), .A1 (nx7367)) ;
    nand02 ix7362 (.Y (nx7361), .A0 (nx2018), .A1 (nx2044)) ;
    nand02 ix2045 (.Y (nx2044), .A0 (nx7365), .A1 (nx7519)) ;
    dffr i5_MR_reg_dataout_15 (.Q (i5_MARo_15), .QB (nx7356), .D (nx2052), .CLK (
         CLK), .R (Rst)) ;
    oai21 ix7371 (.Y (nx7370), .A0 (nx2062), .A1 (nx2060), .B0 (nx7885)) ;
    nor02_2x ix2063 (.Y (nx2062), .A0 (nx7354), .A1 (nx7901)) ;
    nor02_2x ix2061 (.Y (nx2060), .A0 (nx7356), .A1 (nx1642)) ;
    nor02_2x ix7551 (.Y (readenable), .A0 (nx7377), .A1 (nx3563)) ;
    inv01 ix7378 (.Y (nx7377), .A (OuterRead)) ;
    nand02 ix1167 (.Y (EnableReadingFromCPU), .A0 (nx7381), .A1 (nx7383)) ;
    nand03 ix7382 (.Y (nx7381), .A0 (nx7392), .A1 (nx7763), .A2 (nx7907)) ;
    nand03 ix7384 (.Y (nx7383), .A0 (nx7397), .A1 (CNNIMGLOAD), .A2 (nx7907)) ;
    inv02 ix7389 (.Y (nx7390), .A (nx4203)) ;
    inv02 ix7391 (.Y (nx7392), .A (nx4203)) ;
    inv02 ix7393 (.Y (nx7395), .A (nx4083)) ;
    inv02 ix7396 (.Y (nx7397), .A (nx4083)) ;
    inv04 ix7400 (.Y (nx7401), .A (nx7399)) ;
    inv04 ix7402 (.Y (nx7403), .A (nx9396)) ;
    inv04 ix7404 (.Y (nx7405), .A (nx9396)) ;
    inv04 ix7406 (.Y (nx7407), .A (nx9396)) ;
    inv04 ix7408 (.Y (nx7409), .A (nx9396)) ;
    inv04 ix7410 (.Y (nx7411), .A (nx9396)) ;
    inv02 ix7412 (.Y (nx7413), .A (nx7771)) ;
    inv02 ix7414 (.Y (nx7415), .A (nx7771)) ;
    inv01 ix7416 (.Y (nx7417), .A (nx370)) ;
    inv02 ix7418 (.Y (nx7419), .A (nx7417)) ;
    inv02 ix7420 (.Y (nx7421), .A (nx7417)) ;
    inv02 ix7422 (.Y (nx7423), .A (nx7417)) ;
    inv02 ix7424 (.Y (nx7425), .A (nx7417)) ;
    buf02 ix7426 (.Y (nx7427), .A (nx374)) ;
    buf02 ix7428 (.Y (nx7429), .A (nx374)) ;
    buf02 ix7430 (.Y (nx7431), .A (nx374)) ;
    inv02 ix7434 (.Y (nx7435), .A (nx7433)) ;
    inv02 ix7436 (.Y (nx7437), .A (nx7433)) ;
    inv02 ix7438 (.Y (nx7439), .A (nx7433)) ;
    inv02 ix7440 (.Y (nx7441), .A (nx4217)) ;
    inv02 ix7442 (.Y (nx7443), .A (nx4217)) ;
    inv02 ix7444 (.Y (nx7445), .A (nx4217)) ;
    inv02 ix7446 (.Y (nx7447), .A (nx4301)) ;
    inv02 ix7448 (.Y (nx7449), .A (nx4301)) ;
    nand02 ix7450 (.Y (nx7451), .A0 (nx5209), .A1 (nx7857)) ;
    nor02_2x ix7454 (.Y (nx7455), .A0 (nx4532), .A1 (nx7789)) ;
    nor02_2x ix7456 (.Y (nx7457), .A0 (nx4532), .A1 (nx7789)) ;
    nor02_2x ix7458 (.Y (nx7459), .A0 (nx4547), .A1 (nx7789)) ;
    nor02_2x ix7460 (.Y (nx7461), .A0 (nx4547), .A1 (nx7789)) ;
    nor02_2x ix7462 (.Y (nx7463), .A0 (nx4553), .A1 (nx7789)) ;
    nor02_2x ix7464 (.Y (nx7465), .A0 (nx4553), .A1 (nx7791)) ;
    nor02_2x ix7466 (.Y (nx7467), .A0 (nx4558), .A1 (nx7791)) ;
    nor02_2x ix7468 (.Y (nx7469), .A0 (nx4558), .A1 (nx7791)) ;
    nor02_2x ix7470 (.Y (nx7471), .A0 (nx4565), .A1 (nx7791)) ;
    nor02_2x ix7472 (.Y (nx7473), .A0 (nx4565), .A1 (nx7791)) ;
    nor02_2x ix7474 (.Y (nx7475), .A0 (nx4570), .A1 (nx7791)) ;
    nor02_2x ix7476 (.Y (nx7477), .A0 (nx4570), .A1 (nx7791)) ;
    nor02_2x ix7478 (.Y (nx7479), .A0 (nx4577), .A1 (nx7793)) ;
    nor02_2x ix7480 (.Y (nx7481), .A0 (nx4577), .A1 (nx7793)) ;
    nor02_2x ix7482 (.Y (nx7483), .A0 (nx4582), .A1 (nx7793)) ;
    nor02_2x ix7484 (.Y (nx7485), .A0 (nx4582), .A1 (nx7793)) ;
    nor02_2x ix7486 (.Y (nx7487), .A0 (nx4511), .A1 (nx7793)) ;
    nor02_2x ix7488 (.Y (nx7489), .A0 (nx4511), .A1 (nx7793)) ;
    nor02_2x ix7490 (.Y (nx7491), .A0 (nx4592), .A1 (nx7793)) ;
    nor02_2x ix7492 (.Y (nx7493), .A0 (nx4592), .A1 (nx7795)) ;
    nor02_2x ix7494 (.Y (nx7495), .A0 (nx4397), .A1 (nx7795)) ;
    nor02_2x ix7496 (.Y (nx7497), .A0 (nx4397), .A1 (nx7795)) ;
    nor02_2x ix7498 (.Y (nx7499), .A0 (nx4377), .A1 (nx7795)) ;
    nor02_2x ix7500 (.Y (nx7501), .A0 (nx4377), .A1 (nx7795)) ;
    nor02_2x ix7502 (.Y (nx7503), .A0 (nx4381), .A1 (nx7795)) ;
    nor02_2x ix7504 (.Y (nx7505), .A0 (nx4381), .A1 (nx7795)) ;
    nor02_2x ix7506 (.Y (nx7507), .A0 (nx4460), .A1 (nx7797)) ;
    nor02_2x ix7508 (.Y (nx7509), .A0 (nx4460), .A1 (nx7797)) ;
    inv02 ix7510 (.Y (nx7511), .A (nx5259)) ;
    inv02 ix7514 (.Y (nx7515), .A (nx7885)) ;
    inv02 ix7516 (.Y (nx7517), .A (nx7885)) ;
    inv02 ix7518 (.Y (nx7519), .A (nx7885)) ;
    nor02_2x ix7520 (.Y (nx7521), .A0 (nx7095), .A1 (nx7909)) ;
    nor02_2x ix7522 (.Y (nx7523), .A0 (nx7095), .A1 (nx7909)) ;
    buf02 ix7524 (.Y (nx7525), .A (nx1794)) ;
    buf02 ix7526 (.Y (nx7527), .A (nx1906)) ;
    buf02 ix7528 (.Y (nx7529), .A (nx2068)) ;
    buf02 ix7530 (.Y (nx7531), .A (nx2068)) ;
    nand02 ix7536 (.Y (nx7537), .A0 (nx4522), .A1 (nx7857)) ;
    inv01 ix7538 (.Y (nx7539), .A (nx2118)) ;
    inv01 ix7540 (.Y (nx7541), .A (nx7539)) ;
    inv01 ix7550 (.Y (nx7551), .A (nx2238)) ;
    inv02 ix7552 (.Y (nx7553), .A (nx7551)) ;
    inv02 ix7554 (.Y (nx7555), .A (nx7551)) ;
    inv01 ix7556 (.Y (nx7557), .A (nx2264)) ;
    inv02 ix7558 (.Y (nx7559), .A (nx7557)) ;
    inv02 ix7560 (.Y (nx7561), .A (nx7557)) ;
    inv01 ix7562 (.Y (nx7563), .A (nx2290)) ;
    inv02 ix7564 (.Y (nx7565), .A (nx7563)) ;
    inv02 ix7566 (.Y (nx7567), .A (nx7563)) ;
    inv01 ix7568 (.Y (nx7569), .A (nx2320)) ;
    inv01 ix7570 (.Y (nx7571), .A (nx7569)) ;
    nand02 ix7574 (.Y (nx7575), .A0 (nx4613), .A1 (nx7857)) ;
    inv01 ix7576 (.Y (nx7577), .A (nx2520)) ;
    inv01 ix7578 (.Y (nx7579), .A (nx7577)) ;
    inv01 ix7580 (.Y (nx7581), .A (nx2708)) ;
    inv01 ix7582 (.Y (nx7583), .A (nx7581)) ;
    nand02 ix7586 (.Y (nx7587), .A0 (nx4663), .A1 (nx7857)) ;
    inv01 ix7588 (.Y (nx7589), .A (nx2910)) ;
    inv01 ix7590 (.Y (nx7591), .A (nx7589)) ;
    inv01 ix7592 (.Y (nx7593), .A (nx3098)) ;
    inv01 ix7594 (.Y (nx7595), .A (nx7593)) ;
    nand02 ix7598 (.Y (nx7599), .A0 (nx4711), .A1 (nx7857)) ;
    inv01 ix7600 (.Y (nx7601), .A (nx3298)) ;
    inv01 ix7602 (.Y (nx7603), .A (nx7601)) ;
    inv01 ix7604 (.Y (nx7605), .A (nx3486)) ;
    inv01 ix7606 (.Y (nx7607), .A (nx7605)) ;
    nand02 ix7610 (.Y (nx7611), .A0 (nx4757), .A1 (nx7857)) ;
    inv01 ix7612 (.Y (nx7613), .A (nx3698)) ;
    inv01 ix7614 (.Y (nx7615), .A (nx7613)) ;
    inv01 ix7616 (.Y (nx7617), .A (nx3886)) ;
    inv01 ix7618 (.Y (nx7619), .A (nx7617)) ;
    nand02 ix7622 (.Y (nx7623), .A0 (nx4804), .A1 (nx7859)) ;
    inv01 ix7624 (.Y (nx7625), .A (nx4082)) ;
    inv01 ix7626 (.Y (nx7627), .A (nx7625)) ;
    inv01 ix7628 (.Y (nx7629), .A (nx4270)) ;
    inv01 ix7630 (.Y (nx7631), .A (nx7629)) ;
    inv01 ix7634 (.Y (nx7635), .A (nx7633)) ;
    inv01 ix7636 (.Y (nx7637), .A (nx7633)) ;
    inv01 ix7638 (.Y (nx7639), .A (nx7633)) ;
    nand02 ix7642 (.Y (nx7643), .A0 (nx4847), .A1 (nx7859)) ;
    inv01 ix7644 (.Y (nx7645), .A (nx4476)) ;
    inv01 ix7646 (.Y (nx7647), .A (nx7645)) ;
    inv01 ix7648 (.Y (nx7649), .A (nx4664)) ;
    inv01 ix7650 (.Y (nx7651), .A (nx7649)) ;
    nand02 ix7654 (.Y (nx7655), .A0 (nx4894), .A1 (nx7859)) ;
    inv01 ix7656 (.Y (nx7657), .A (nx4860)) ;
    inv01 ix7658 (.Y (nx7659), .A (nx7657)) ;
    inv01 ix7660 (.Y (nx7661), .A (nx5048)) ;
    inv01 ix7662 (.Y (nx7663), .A (nx7661)) ;
    nand02 ix7666 (.Y (nx7667), .A0 (nx4937), .A1 (nx7859)) ;
    inv01 ix7668 (.Y (nx7669), .A (nx5258)) ;
    inv01 ix7670 (.Y (nx7671), .A (nx7669)) ;
    inv01 ix7672 (.Y (nx7673), .A (nx5446)) ;
    inv01 ix7674 (.Y (nx7675), .A (nx7673)) ;
    nand02 ix7678 (.Y (nx7679), .A0 (nx4985), .A1 (nx7859)) ;
    inv01 ix7680 (.Y (nx7681), .A (nx5642)) ;
    inv01 ix7682 (.Y (nx7683), .A (nx7681)) ;
    inv01 ix7684 (.Y (nx7685), .A (nx5830)) ;
    inv01 ix7686 (.Y (nx7687), .A (nx7685)) ;
    nand02 ix7690 (.Y (nx7691), .A0 (nx5029), .A1 (nx7859)) ;
    inv01 ix7692 (.Y (nx7693), .A (nx6032)) ;
    inv01 ix7694 (.Y (nx7695), .A (nx7693)) ;
    inv01 ix7696 (.Y (nx7697), .A (nx6220)) ;
    inv01 ix7698 (.Y (nx7699), .A (nx7697)) ;
    nand02 ix7702 (.Y (nx7703), .A0 (nx5075), .A1 (nx7859)) ;
    inv01 ix7704 (.Y (nx7705), .A (nx6416)) ;
    inv01 ix7706 (.Y (nx7707), .A (nx7705)) ;
    inv01 ix7708 (.Y (nx7709), .A (nx6604)) ;
    inv01 ix7710 (.Y (nx7711), .A (nx7709)) ;
    nand02 ix7714 (.Y (nx7715), .A0 (nx5119), .A1 (nx7861)) ;
    inv01 ix7716 (.Y (nx7717), .A (nx6808)) ;
    inv01 ix7718 (.Y (nx7719), .A (nx7717)) ;
    inv01 ix7720 (.Y (nx7721), .A (nx6996)) ;
    inv01 ix7722 (.Y (nx7723), .A (nx7721)) ;
    nand02 ix7726 (.Y (nx7727), .A0 (nx5165), .A1 (nx7861)) ;
    inv01 ix7728 (.Y (nx7729), .A (nx7192)) ;
    inv01 ix7730 (.Y (nx7731), .A (nx7729)) ;
    inv01 ix7732 (.Y (nx7733), .A (nx7380)) ;
    inv01 ix7734 (.Y (nx7735), .A (nx7733)) ;
    buf02 ix7736 (.Y (nx7737), .A (nx3523)) ;
    buf02 ix7738 (.Y (nx7739), .A (nx3523)) ;
    inv02 ix7740 (.Y (nx7741), .A (CNNIMGLOAD)) ;
    inv02 ix7742 (.Y (nx7743), .A (CNNIMGLOAD)) ;
    inv02 ix7744 (.Y (nx7745), .A (CNNIMGLOAD)) ;
    inv02 ix7746 (.Y (nx7747), .A (CNNIMGLOAD)) ;
    inv02 ix7748 (.Y (nx7749), .A (CNNIMGLOAD)) ;
    inv02 ix7750 (.Y (nx7751), .A (CNNIMGLOAD)) ;
    inv02 ix7752 (.Y (nx7753), .A (CNNIMGLOAD)) ;
    inv02 ix7754 (.Y (nx7755), .A (CNNIMGLOAD)) ;
    inv02 ix7756 (.Y (nx7757), .A (CNNIMGLOAD)) ;
    inv02 ix7758 (.Y (nx7759), .A (CNNIMGLOAD)) ;
    inv02 ix7760 (.Y (nx7761), .A (CNNIMGLOAD)) ;
    inv02 ix7762 (.Y (nx7763), .A (CNNIMGLOAD)) ;
    nor02_2x ix7764 (.Y (nx7765), .A0 (nx3093), .A1 (nx282)) ;
    nor02_2x ix7766 (.Y (nx7767), .A0 (nx3093), .A1 (nx282)) ;
    inv02 ix7768 (.Y (nx7769), .A (i8_reset1)) ;
    inv02 ix7770 (.Y (nx7771), .A (i8_reset1)) ;
    inv01 ix7772 (.Y (nx7773), .A (nx3921)) ;
    inv02 ix7774 (.Y (nx7775), .A (nx7773)) ;
    inv02 ix7776 (.Y (nx7777), .A (nx7773)) ;
    inv02 ix7778 (.Y (nx7779), .A (nx7773)) ;
    nor02_2x ix7780 (.Y (nx7781), .A0 (nx3940), .A1 (nx4126)) ;
    inv02 ix7784 (.Y (nx7785), .A (nx7783)) ;
    inv02 ix7786 (.Y (nx7787), .A (nx7783)) ;
    inv02 ix7788 (.Y (nx7789), .A (nx7783)) ;
    inv02 ix7790 (.Y (nx7791), .A (nx7783)) ;
    inv02 ix7792 (.Y (nx7793), .A (nx7783)) ;
    inv02 ix7794 (.Y (nx7795), .A (nx7783)) ;
    inv02 ix7796 (.Y (nx7797), .A (nx7783)) ;
    buf02 ix7798 (.Y (nx7799), .A (nx3971)) ;
    buf02 ix7800 (.Y (nx7801), .A (nx3971)) ;
    buf02 ix7802 (.Y (nx7803), .A (nx3999)) ;
    buf02 ix7804 (.Y (nx7805), .A (nx3999)) ;
    inv02 ix7806 (.Y (nx7807), .A (i8_counterout2_2)) ;
    inv02 ix7808 (.Y (nx7809), .A (nx7913)) ;
    nand02 ix7810 (.Y (nx7811), .A0 (i8_reset2), .A1 (zed)) ;
    nor02_2x ix7812 (.Y (nx7813), .A0 (i8_counterout2_0), .A1 (i8_counterout2_1)
             ) ;
    inv02 ix7814 (.Y (nx7815), .A (i8_counterout2_3)) ;
    inv02 ix7816 (.Y (nx7817), .A (i8_counterout2_3)) ;
    inv02 ix7818 (.Y (nx7819), .A (i7_start)) ;
    inv02 ix7820 (.Y (nx7821), .A (i7_start)) ;
    inv02 ix7822 (.Y (nx7823), .A (i7_start)) ;
    buf02 ix7824 (.Y (nx7825), .A (nx4246)) ;
    buf02 ix7826 (.Y (nx7827), .A (nx4246)) ;
    buf02 ix7828 (.Y (nx7829), .A (nx4271)) ;
    buf02 ix7830 (.Y (nx7831), .A (nx4271)) ;
    buf02 ix7832 (.Y (nx7833), .A (nx4274)) ;
    buf02 ix7834 (.Y (nx7835), .A (nx4274)) ;
    nor02_2x ix7836 (.Y (nx7837), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)
             ) ;
    buf02 ix7838 (.Y (nx7839), .A (nx4303)) ;
    buf02 ix7840 (.Y (nx7841), .A (nx4303)) ;
    buf02 ix7842 (.Y (nx7843), .A (nx4405)) ;
    buf02 ix7844 (.Y (nx7845), .A (nx4405)) ;
    buf02 ix7846 (.Y (nx7847), .A (nx4407)) ;
    buf02 ix7848 (.Y (nx7849), .A (nx4407)) ;
    inv02 ix7852 (.Y (nx7853), .A (nx7851)) ;
    inv02 ix7854 (.Y (nx7855), .A (nx7851)) ;
    inv02 ix7856 (.Y (nx7857), .A (nx7851)) ;
    inv02 ix7858 (.Y (nx7859), .A (nx7851)) ;
    inv02 ix7860 (.Y (nx7861), .A (nx7851)) ;
    nor02_2x ix7862 (.Y (nx7863), .A0 (nx3940), .A1 (i8_counterout2_1)) ;
    nor02_2x ix7864 (.Y (nx7865), .A0 (i8_counterout2_0), .A1 (nx4126)) ;
    inv02 ix7868 (.Y (nx7869), .A (nx7867)) ;
    inv02 ix7870 (.Y (nx7871), .A (nx7867)) ;
    inv02 ix7872 (.Y (nx7873), .A (nx7867)) ;
    inv02 ix7874 (.Y (nx7875), .A (nx7867)) ;
    inv02 ix7876 (.Y (nx7877), .A (i5_FAEN)) ;
    inv02 ix7878 (.Y (nx7879), .A (i5_FAEN)) ;
    inv02 ix7880 (.Y (nx7881), .A (i5_FAEN)) ;
    inv02 ix7882 (.Y (nx7883), .A (i5_FAEN)) ;
    inv02 ix7884 (.Y (nx7885), .A (i5_FAEN)) ;
    inv02 ix7888 (.Y (nx7889), .A (nx7887)) ;
    inv02 ix7890 (.Y (nx7891), .A (nx9398)) ;
    inv02 ix7892 (.Y (nx7893), .A (nx9398)) ;
    inv02 ix7894 (.Y (nx7895), .A (nx9398)) ;
    inv02 ix7896 (.Y (nx7897), .A (nx9398)) ;
    inv02 ix7898 (.Y (nx7899), .A (nx9398)) ;
    inv02 ix7900 (.Y (nx7901), .A (nx9398)) ;
    inv02 ix7906 (.Y (nx7907), .A (nx7959)) ;
    inv02 ix7908 (.Y (nx7909), .A (nx7959)) ;
    inv02 ix7910 (.Y (nx7911), .A (nx7807)) ;
    inv02 ix7912 (.Y (nx7913), .A (nx7807)) ;
    inv02 ix7956 (.Y (nx7957), .A (loadenable)) ;
    inv02 ix7958 (.Y (nx7959), .A (loadenable)) ;
    inv02 ix7960 (.Y (nx7961), .A (i8_counterout2_2)) ;
    nor02_2x ix3524 (.Y (nx3523), .A0 (nx66), .A1 (Rst)) ;
    nor02_2x ix69 (.Y (nx7399), .A0 (nx8009), .A1 (Rst)) ;
    inv01 ix8008 (.Y (nx8009), .A (nx3565)) ;
    nor02_2x ix3936 (.Y (nx3935), .A0 (nx528), .A1 (nx4151)) ;
    nor02_2x ix3944 (.Y (nx3943), .A0 (nx376), .A1 (nx3940)) ;
    nand02 ix3953 (.Y (nx7783), .A0 (nx8011), .A1 (nx7779)) ;
    aoi21 ix369 (.Y (nx8011), .A0 (i8_reset2), .A1 (zed), .B0 (nx4083)) ;
    mux21 ix3158 (.Y (nx3157), .A0 (nx8013), .A1 (nx3967), .S0 (nx7803)) ;
    inv01 ix8012 (.Y (nx8013), .A (nx206)) ;
    mux21 ix3178 (.Y (nx3177), .A0 (nx8015), .A1 (nx3979), .S0 (nx7803)) ;
    inv01 ix8014 (.Y (nx8015), .A (nx254)) ;
    nor02_2x ix4014 (.Y (nx4013), .A0 (nx3092), .A1 (i8_counterout1_3)) ;
    nor02_2x ix4030 (.Y (nx4029), .A0 (nx314), .A1 (nx7773)) ;
    mux21 ix3148 (.Y (nx3147), .A0 (nx8017), .A1 (nx4033), .S0 (nx7803)) ;
    inv01 ix8016 (.Y (nx8017), .A (nx182)) ;
    mux21 ix3168 (.Y (nx3167), .A0 (nx8019), .A1 (nx4050), .S0 (nx7803)) ;
    inv01 ix8018 (.Y (nx8019), .A (nx230)) ;
    xnor2 ix4067 (.Y (nx4066), .A0 (nx4059), .A1 (nx8021)) ;
    nand02 ix4070 (.Y (nx8021), .A0 (nx8023), .A1 (nx3979)) ;
    inv01 ix8022 (.Y (nx8023), .A (nx3097)) ;
    nor02_2x ix4080 (.Y (nx4079), .A0 (nx3095), .A1 (i8_counterout1_5)) ;
    xnor2 ix397 (.Y (nx396), .A0 (nx3940), .A1 (nx4126)) ;
    xnor2 ix445 (.Y (nx444), .A0 (nx4151), .A1 (nx8025)) ;
    inv01 ix8024 (.Y (nx8025), .A (nx3101)) ;
    xnor2 ix481 (.Y (nx480), .A0 (nx4167), .A1 (nx8027)) ;
    inv01 ix8026 (.Y (nx8027), .A (nx458)) ;
    xnor2 ix465 (.Y (nx464), .A0 (nx4159), .A1 (nx8029)) ;
    inv01 ix8028 (.Y (nx8029), .A (nx3100)) ;
    xnor2 ix495 (.Y (nx494), .A0 (nx4177), .A1 (nx8031)) ;
    nor02_2x ix493 (.Y (nx8031), .A0 (nx8033), .A1 (i8_counterout2_6)) ;
    nand02 ix4176 (.Y (nx8033), .A0 (nx8029), .A1 (nx4159)) ;
    nor02_2x ix4199 (.Y (nx4198), .A0 (nx602), .A1 (nx7773)) ;
    xnor2 ix725 (.Y (nx724), .A0 (nx4283), .A1 (nx8035)) ;
    inv01 ix8034 (.Y (nx8035), .A (nx3111)) ;
    nor02_2x ix4299 (.Y (nx4298), .A0 (nx654), .A1 (nx4309)) ;
    nor02_2x ix4304 (.Y (nx4303), .A0 (nx648), .A1 (i7_start)) ;
    xnor2 ix675 (.Y (nx674), .A0 (nx4309), .A1 (nx4317)) ;
    xnor2 ix709 (.Y (nx708), .A0 (nx4318), .A1 (nx8037)) ;
    nor03_2x ix703 (.Y (nx8037), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)
             , .A2 (i7_counterout2_2)) ;
    xnor2 ix741 (.Y (nx740), .A0 (nx4333), .A1 (nx8039)) ;
    inv01 ix8038 (.Y (nx8039), .A (nx3109)) ;
    xnor2 ix759 (.Y (nx758), .A0 (nx4345), .A1 (nx8041)) ;
    inv01 ix8040 (.Y (nx8041), .A (nx3107)) ;
    xnor2 ix773 (.Y (nx772), .A0 (nx4355), .A1 (nx8043)) ;
    nor02_2x ix771 (.Y (nx8043), .A0 (nx8045), .A1 (i7_counterout2_6)) ;
    nand02 ix4366 (.Y (nx8045), .A0 (nx8039), .A1 (nx4333)) ;
    nand03 ix897 (.Y (nx4383), .A0 (DataBus[12]), .A1 (DataBus[11]), .A2 (nx8047
           )) ;
    inv01 ix8046 (.Y (nx8047), .A (nx4379)) ;
    nor02_2x ix4387 (.Y (nx4386), .A0 (nx3117), .A1 (i7_counterout1_4)) ;
    nor02_2x ix4408 (.Y (nx4407), .A0 (nx856), .A1 (i7_start)) ;
    nor02_2x ix4420 (.Y (nx4419), .A0 (nx3118), .A1 (i7_counterout1_3)) ;
    nor02_2x ix4438 (.Y (nx4437), .A0 (nx3116), .A1 (i7_counterout1_5)) ;
    nor02_2x ix4463 (.Y (nx4462), .A0 (nx3115), .A1 (i7_counterout1_6)) ;
    xnor2 ix1101 (.Y (nx1100), .A0 (nx4487), .A1 (nx8049)) ;
    nor02_2x ix1099 (.Y (nx8049), .A0 (nx8051), .A1 (i7_counterout1_6)) ;
    inv01 ix8050 (.Y (nx8051), .A (nx4437)) ;
    xnor2 ix691 (.Y (nx690), .A0 (nx4239), .A1 (nx8053)) ;
    nor02_2x ix685 (.Y (nx8053), .A0 (i7_counterout2_0), .A1 (i7_counterout2_1)
             ) ;
    nand03 ix551 (.Y (nx7433), .A0 (nx4191), .A1 (nx8055), .A2 (
           EnableReadingFromCPU2)) ;
    inv01 ix8054 (.Y (nx8055), .A (DataBus[15])) ;
    nand03 ix4530 (.Y (nx7851), .A0 (nx3925), .A1 (CNNIMGLOAD), .A2 (nx9396)) ;
    nor02_2x ix1399 (.Y (nx1398), .A0 (nx7511), .A1 (nx8057)) ;
    inv01 ix8056 (.Y (nx8057), .A (nx1188)) ;
    nor02_2x ix1411 (.Y (nx1410), .A0 (nx7511), .A1 (nx8059)) ;
    inv01 ix8058 (.Y (nx8059), .A (nx1202)) ;
    nor02_2x ix1423 (.Y (nx1422), .A0 (nx7511), .A1 (nx8061)) ;
    inv01 ix8060 (.Y (nx8061), .A (nx1216)) ;
    nor02_2x ix1435 (.Y (nx1434), .A0 (nx7511), .A1 (nx8063)) ;
    inv01 ix8062 (.Y (nx8063), .A (nx1230)) ;
    nor02_2x ix1447 (.Y (nx1446), .A0 (nx7511), .A1 (nx8065)) ;
    inv01 ix8064 (.Y (nx8065), .A (nx1244)) ;
    nor02_2x ix1459 (.Y (nx1458), .A0 (nx7511), .A1 (nx8067)) ;
    inv01 ix8066 (.Y (nx8067), .A (nx1258)) ;
    nor02_2x ix1471 (.Y (nx1470), .A0 (nx7511), .A1 (nx8069)) ;
    inv01 ix8068 (.Y (nx8069), .A (nx1272)) ;
    nor02_2x ix1483 (.Y (nx1482), .A0 (nx1388), .A1 (nx8071)) ;
    inv01 ix8070 (.Y (nx8071), .A (nx1286)) ;
    nor02_2x ix1495 (.Y (nx1494), .A0 (nx1388), .A1 (nx8073)) ;
    inv01 ix8072 (.Y (nx8073), .A (nx1300)) ;
    nor02_2x ix1507 (.Y (nx1506), .A0 (nx1388), .A1 (nx8075)) ;
    inv01 ix8074 (.Y (nx8075), .A (nx1314)) ;
    nor02_2x ix1519 (.Y (nx1518), .A0 (nx1388), .A1 (nx8077)) ;
    inv01 ix8076 (.Y (nx8077), .A (nx1328)) ;
    nor02_2x ix1531 (.Y (nx1530), .A0 (nx1388), .A1 (nx8079)) ;
    inv01 ix8078 (.Y (nx8079), .A (nx1342)) ;
    nor02_2x ix1543 (.Y (nx1542), .A0 (nx1388), .A1 (nx8081)) ;
    inv01 ix8080 (.Y (nx8081), .A (nx1356)) ;
    nor02_2x ix1555 (.Y (nx1554), .A0 (nx1388), .A1 (nx8083)) ;
    inv01 ix8082 (.Y (nx8083), .A (nx1370)) ;
    nand03 ix5312 (.Y (nx7867), .A0 (nx4227), .A1 (nx7741), .A2 (nx9396)) ;
    nand03 ix4445 (.Y (nx7633), .A0 (nx8085), .A1 (nx4283), .A2 (nx8087)) ;
    inv01 ix8084 (.Y (nx8085), .A (nx7845)) ;
    inv01 ix8086 (.Y (nx8087), .A (nx7841)) ;
    mux21 ix1651 (.Y (Address[0]), .A0 (nx7039), .A1 (nx7037), .S0 (nx9398)) ;
    xnor2 ix1635 (.Y (nx1634), .A0 (nx7885), .A1 (nx8089)) ;
    inv01 ix8088 (.Y (nx8089), .A (nx7072)) ;
    nor02_2x ix7056 (.Y (NOT_nx814), .A0 (nx812), .A1 (i7_tmp)) ;
    mux21 ix7073 (.Y (nx7072), .A0 (i5_MARo_0), .A1 (OuterAddress[0]), .S0 (
          nx9400)) ;
    nor02_2x ix7076 (.Y (nx7887), .A0 (nx7095), .A1 (loadenable)) ;
    mux21 ix1673 (.Y (Address[1]), .A0 (nx7081), .A1 (nx7079), .S0 (nx9400)) ;
    mux21 ix1701 (.Y (Address[2]), .A0 (nx7100), .A1 (nx7098), .S0 (nx9400)) ;
    mux21 ix7108 (.Y (nx7107), .A0 (i5_MARo_1), .A1 (OuterAddress[1]), .S0 (
          nx9400)) ;
    mux21 ix1729 (.Y (Address[3]), .A0 (nx7117), .A1 (nx7115), .S0 (nx9400)) ;
    mux21 ix7127 (.Y (nx7126), .A0 (i5_MARo_2), .A1 (OuterAddress[2]), .S0 (
          nx9400)) ;
    mux21 ix7130 (.Y (nx7129), .A0 (i5_MARo_3), .A1 (OuterAddress[3]), .S0 (
          nx9400)) ;
    mux21 ix1757 (.Y (Address[4]), .A0 (nx7139), .A1 (nx7137), .S0 (nx9402)) ;
    mux21 ix7149 (.Y (nx7148), .A0 (i5_MARo_4), .A1 (OuterAddress[4]), .S0 (
          nx9402)) ;
    mux21 ix1785 (.Y (Address[5]), .A0 (nx7159), .A1 (nx7157), .S0 (nx9402)) ;
    mux21 ix7170 (.Y (nx7169), .A0 (i5_MARo_5), .A1 (OuterAddress[5]), .S0 (
          nx9402)) ;
    mux21 ix1813 (.Y (Address[6]), .A0 (nx7181), .A1 (nx7178), .S0 (nx9402)) ;
    mux21 ix1841 (.Y (Address[7]), .A0 (nx7199), .A1 (nx7197), .S0 (nx9402)) ;
    mux21 ix7210 (.Y (nx7209), .A0 (i5_MARo_6), .A1 (OuterAddress[6]), .S0 (
          nx9402)) ;
    mux21 ix7212 (.Y (nx7211), .A0 (i5_MARo_7), .A1 (OuterAddress[7]), .S0 (
          nx9404)) ;
    mux21 ix1869 (.Y (Address[8]), .A0 (nx7223), .A1 (nx7221), .S0 (nx9404)) ;
    mux21 ix7234 (.Y (nx7233), .A0 (i5_MARo_8), .A1 (OuterAddress[8]), .S0 (
          nx9404)) ;
    mux21 ix1897 (.Y (Address[9]), .A0 (nx7243), .A1 (nx7241), .S0 (nx9404)) ;
    mux21 ix7254 (.Y (nx7253), .A0 (i5_MARo_9), .A1 (OuterAddress[9]), .S0 (
          nx9404)) ;
    mux21 ix1925 (.Y (Address[10]), .A0 (nx7265), .A1 (nx7262), .S0 (nx9404)) ;
    mux21 ix1953 (.Y (Address[11]), .A0 (nx7279), .A1 (nx7277), .S0 (nx9404)) ;
    mux21 ix7288 (.Y (nx7287), .A0 (i5_MARo_10), .A1 (OuterAddress[10]), .S0 (
          nx9406)) ;
    mux21 ix7290 (.Y (nx7289), .A0 (i5_MARo_11), .A1 (OuterAddress[11]), .S0 (
          nx9406)) ;
    mux21 ix1981 (.Y (Address[12]), .A0 (nx7301), .A1 (nx7298), .S0 (nx9406)) ;
    mux21 ix7311 (.Y (nx7310), .A0 (i5_MARo_12), .A1 (OuterAddress[12]), .S0 (
          nx9406)) ;
    mux21 ix2009 (.Y (Address[13]), .A0 (nx7321), .A1 (nx7319), .S0 (nx9406)) ;
    mux21 ix7331 (.Y (nx7330), .A0 (i5_MARo_13), .A1 (OuterAddress[13]), .S0 (
          nx9406)) ;
    mux21 ix2037 (.Y (Address[14]), .A0 (nx7341), .A1 (nx7339), .S0 (nx9406)) ;
    mux21 ix2065 (.Y (Address[15]), .A0 (nx7356), .A1 (nx7354), .S0 (nx9408)) ;
    mux21 ix7366 (.Y (nx7365), .A0 (i5_MARo_14), .A1 (OuterAddress[14]), .S0 (
          nx9408)) ;
    mux21 ix7368 (.Y (nx7367), .A0 (i5_MARo_15), .A1 (OuterAddress[15]), .S0 (
          nx9408)) ;
    latchr i8_lat_reset1_u1 (.QB (nx5), .D (i8_nx74), .CLK (nx298), .R (
           DecompressedData1[255])) ;
    inv01 i8_lat_reset1_u2 (.Y (i8_reset1), .A (nx5)) ;
    latchs_ni i8_lat_tmp_u1 (.QB (nx8093), .D (DecompressedData1[255]), .CLK (
              nx536), .S (nx540)) ;
    inv02 i8_lat_tmp_u2 (.Y (zed), .A (nx8093)) ;
    buf02 i8_lat_tmp_u3 (.Y (nx3955), .A (nx8093)) ;
    latchs_ni i7_lat_tmp_u1 (.QB (nx8096), .D (DecompressedData1[255]), .CLK (
              nx1140), .S (nx1148)) ;
    inv02 i7_lat_tmp_u2 (.Y (i7_tmp), .A (nx8096)) ;
    buf02 i7_lat_tmp_u3 (.Y (nx4277), .A (nx8096)) ;
    latchr i7_r28_lat_q_0__u1 (.QB (nx8099), .D (nx9280), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_0__u2 (.Y (DecompressedData1[0]), .A (nx8099)) ;
    buf02 i7_r28_lat_q_0__u3 (.Y (nx5695), .A (nx8099)) ;
    latchr i8_r1_lat_q_0__u1 (.QB (nx8102), .D (nx2122), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_0__u2 (.Y (DecompressedData2[0]), .A (nx8102)) ;
    buf02 i8_r1_lat_q_0__u3 (.Y (nx5697), .A (nx8102)) ;
    latchr i7_r28_lat_q_1__u1 (.QB (nx8105), .D (nx9294), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_1__u2 (.Y (DecompressedData1[1]), .A (nx8105)) ;
    buf02 i7_r28_lat_q_1__u3 (.Y (nx5700), .A (nx8105)) ;
    latchr i8_r1_lat_q_1__u1 (.QB (nx8108), .D (nx2148), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_1__u2 (.Y (DecompressedData2[1]), .A (nx8108)) ;
    buf02 i8_r1_lat_q_1__u3 (.Y (nx5703), .A (nx8108)) ;
    latchr i7_r28_lat_q_2__u1 (.QB (nx8111), .D (nx9304), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_2__u2 (.Y (DecompressedData1[2]), .A (nx8111)) ;
    buf02 i7_r28_lat_q_2__u3 (.Y (nx5707), .A (nx8111)) ;
    latchr i8_r1_lat_q_2__u1 (.QB (nx8114), .D (nx2174), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_2__u2 (.Y (DecompressedData2[2]), .A (nx8114)) ;
    buf02 i8_r1_lat_q_2__u3 (.Y (nx5709), .A (nx8114)) ;
    latchr i7_r28_lat_q_3__u1 (.QB (nx8117), .D (nx9314), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_3__u2 (.Y (DecompressedData1[3]), .A (nx8117)) ;
    buf02 i7_r28_lat_q_3__u3 (.Y (nx5712), .A (nx8117)) ;
    latchr i8_r1_lat_q_3__u1 (.QB (nx8120), .D (nx2200), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_3__u2 (.Y (DecompressedData2[3]), .A (nx8120)) ;
    buf02 i8_r1_lat_q_3__u3 (.Y (nx5715), .A (nx8120)) ;
    latchr i7_r28_lat_q_4__u1 (.QB (nx8123), .D (nx9324), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_4__u2 (.Y (DecompressedData1[4]), .A (nx8123)) ;
    buf02 i7_r28_lat_q_4__u3 (.Y (nx5719), .A (nx8123)) ;
    latchr i8_r1_lat_q_4__u1 (.QB (nx8126), .D (nx2226), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_4__u2 (.Y (DecompressedData2[4]), .A (nx8126)) ;
    buf02 i8_r1_lat_q_4__u3 (.Y (nx5721), .A (nx8126)) ;
    latchr i7_r28_lat_q_5__u1 (.QB (nx8129), .D (nx9332), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_5__u2 (.Y (DecompressedData1[5]), .A (nx8129)) ;
    buf02 i7_r28_lat_q_5__u3 (.Y (nx5724), .A (nx8129)) ;
    latchr i8_r1_lat_q_5__u1 (.QB (nx8132), .D (nx2252), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_5__u2 (.Y (DecompressedData2[5]), .A (nx8132)) ;
    buf02 i8_r1_lat_q_5__u3 (.Y (nx5727), .A (nx8132)) ;
    latchr i7_r28_lat_q_6__u1 (.QB (nx8135), .D (nx9336), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_6__u2 (.Y (DecompressedData1[6]), .A (nx8135)) ;
    buf02 i7_r28_lat_q_6__u3 (.Y (nx5731), .A (nx8135)) ;
    latchr i8_r1_lat_q_6__u1 (.QB (nx8138), .D (nx2278), .CLK (nx9288), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_6__u2 (.Y (DecompressedData2[6]), .A (nx8138)) ;
    buf02 i8_r1_lat_q_6__u3 (.Y (nx5733), .A (nx8138)) ;
    latchr i7_r28_lat_q_7__u1 (.QB (nx8141), .D (nx9340), .CLK (nx2080), .R (
           DecompressedData1[255])) ;
    inv01 i7_r28_lat_q_7__u2 (.Y (DecompressedData1[7]), .A (nx8141)) ;
    buf02 i7_r28_lat_q_7__u3 (.Y (nx5736), .A (nx8141)) ;
    latchr i8_r1_lat_q_7__u1 (.QB (nx8144), .D (nx2304), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_7__u2 (.Y (DecompressedData2[7]), .A (nx8144)) ;
    buf02 i8_r1_lat_q_7__u3 (.Y (nx5739), .A (nx8144)) ;
    latchr i7_r27_lat_q_0__u1 (.QB (nx8147), .D (nx9280), .CLK (nx2320), .R (
           DecompressedData1[255])) ;
    inv01 i7_r27_lat_q_0__u2 (.Y (DecompressedData1[8]), .A (nx8147)) ;
    buf02 i7_r27_lat_q_0__u3 (.Y (nx5743), .A (nx8147)) ;
    latchr i8_r1_lat_q_8__u1 (.QB (nx8150), .D (nx2334), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_8__u2 (.Y (DecompressedData2[8]), .A (nx8150)) ;
    buf02 i8_r1_lat_q_8__u3 (.Y (nx5745), .A (nx8150)) ;
    latchr i7_r27_lat_q_1__u1 (.QB (nx8153), .D (nx9294), .CLK (nx2320), .R (
           DecompressedData1[255])) ;
    inv01 i7_r27_lat_q_1__u2 (.Y (DecompressedData1[9]), .A (nx8153)) ;
    buf02 i7_r27_lat_q_1__u3 (.Y (nx5748), .A (nx8153)) ;
    latchr i8_r1_lat_q_9__u1 (.QB (nx8156), .D (nx2358), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_9__u2 (.Y (DecompressedData2[9]), .A (nx8156)) ;
    buf02 i8_r1_lat_q_9__u3 (.Y (nx5751), .A (nx8156)) ;
    latchr i7_r27_lat_q_2__u1 (.QB (nx8159), .D (nx9304), .CLK (nx2320), .R (
           DecompressedData1[255])) ;
    inv01 i7_r27_lat_q_2__u2 (.Y (DecompressedData1[10]), .A (nx8159)) ;
    buf02 i7_r27_lat_q_2__u3 (.Y (nx5755), .A (nx8159)) ;
    latchr i8_r1_lat_q_10__u1 (.QB (nx8162), .D (nx2382), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_10__u2 (.Y (DecompressedData2[10]), .A (nx8162)) ;
    buf02 i8_r1_lat_q_10__u3 (.Y (nx5757), .A (nx8162)) ;
    latchr i7_r27_lat_q_3__u1 (.QB (nx8165), .D (nx9314), .CLK (nx2320), .R (
           DecompressedData1[255])) ;
    inv01 i7_r27_lat_q_3__u2 (.Y (DecompressedData1[11]), .A (nx8165)) ;
    buf02 i7_r27_lat_q_3__u3 (.Y (nx5760), .A (nx8165)) ;
    latchr i8_r1_lat_q_11__u1 (.QB (nx8168), .D (nx2406), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_11__u2 (.Y (DecompressedData2[11]), .A (nx8168)) ;
    buf02 i8_r1_lat_q_11__u3 (.Y (nx5763), .A (nx8168)) ;
    latchr i7_r27_lat_q_4__u1 (.QB (nx8171), .D (nx9324), .CLK (nx2320), .R (
           DecompressedData1[255])) ;
    inv01 i7_r27_lat_q_4__u2 (.Y (DecompressedData1[12]), .A (nx8171)) ;
    buf02 i7_r27_lat_q_4__u3 (.Y (nx5767), .A (nx8171)) ;
    latchr i8_r1_lat_q_12__u1 (.QB (nx8174), .D (nx2430), .CLK (nx9290), .R (
           DecompressedData1[255])) ;
    inv01 i8_r1_lat_q_12__u2 (.Y (DecompressedData2[12]), .A (nx8174)) ;
    buf02 i8_r1_lat_q_12__u3 (.Y (nx5769), .A (nx8174)) ;
    latchr i7_r26_lat_q_0__u1 (.QB (nx8177), .D (nx9280), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_0__u2 (.Y (DecompressedData1[16]), .A (nx8177)) ;
    buf02 i7_r26_lat_q_0__u3 (.Y (nx5785), .A (nx8177)) ;
    latchr i8_r2_lat_q_0__u1 (.QB (nx8180), .D (nx2524), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_0__u2 (.Y (DecompressedData2[16]), .A (nx8180)) ;
    buf02 i8_r2_lat_q_0__u3 (.Y (nx5787), .A (nx8180)) ;
    latchr i7_r26_lat_q_1__u1 (.QB (nx8183), .D (nx9294), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_1__u2 (.Y (DecompressedData1[17]), .A (nx8183)) ;
    buf02 i7_r26_lat_q_1__u3 (.Y (nx5791), .A (nx8183)) ;
    latchr i8_r2_lat_q_1__u1 (.QB (nx8186), .D (nx2548), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_1__u2 (.Y (DecompressedData2[17]), .A (nx8186)) ;
    buf02 i8_r2_lat_q_1__u3 (.Y (nx5793), .A (nx8186)) ;
    latchr i7_r26_lat_q_2__u1 (.QB (nx8189), .D (nx9304), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_2__u2 (.Y (DecompressedData1[18]), .A (nx8189)) ;
    buf02 i7_r26_lat_q_2__u3 (.Y (nx5796), .A (nx8189)) ;
    latchr i8_r2_lat_q_2__u1 (.QB (nx8192), .D (nx2572), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_2__u2 (.Y (DecompressedData2[18]), .A (nx8192)) ;
    buf02 i8_r2_lat_q_2__u3 (.Y (nx5799), .A (nx8192)) ;
    latchr i7_r26_lat_q_3__u1 (.QB (nx8195), .D (nx9314), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_3__u2 (.Y (DecompressedData1[19]), .A (nx8195)) ;
    buf02 i7_r26_lat_q_3__u3 (.Y (nx5803), .A (nx8195)) ;
    latchr i8_r2_lat_q_3__u1 (.QB (nx8198), .D (nx2596), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_3__u2 (.Y (DecompressedData2[19]), .A (nx8198)) ;
    buf02 i8_r2_lat_q_3__u3 (.Y (nx5805), .A (nx8198)) ;
    latchr i7_r26_lat_q_4__u1 (.QB (nx8201), .D (nx9324), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_4__u2 (.Y (DecompressedData1[20]), .A (nx8201)) ;
    buf02 i7_r26_lat_q_4__u3 (.Y (nx5808), .A (nx8201)) ;
    latchr i8_r2_lat_q_4__u1 (.QB (nx8204), .D (nx2620), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_4__u2 (.Y (DecompressedData2[20]), .A (nx8204)) ;
    buf02 i8_r2_lat_q_4__u3 (.Y (nx5811), .A (nx8204)) ;
    latchr i7_r26_lat_q_5__u1 (.QB (nx8207), .D (nx9332), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_5__u2 (.Y (DecompressedData1[21]), .A (nx8207)) ;
    buf02 i7_r26_lat_q_5__u3 (.Y (nx5815), .A (nx8207)) ;
    latchr i8_r2_lat_q_5__u1 (.QB (nx8210), .D (nx2644), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_5__u2 (.Y (DecompressedData2[21]), .A (nx8210)) ;
    buf02 i8_r2_lat_q_5__u3 (.Y (nx5817), .A (nx8210)) ;
    latchr i7_r26_lat_q_6__u1 (.QB (nx8213), .D (nx9336), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_6__u2 (.Y (DecompressedData1[22]), .A (nx8213)) ;
    buf02 i7_r26_lat_q_6__u3 (.Y (nx5820), .A (nx8213)) ;
    latchr i8_r2_lat_q_6__u1 (.QB (nx8216), .D (nx2668), .CLK (nx9344), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_6__u2 (.Y (DecompressedData2[22]), .A (nx8216)) ;
    buf02 i8_r2_lat_q_6__u3 (.Y (nx5823), .A (nx8216)) ;
    latchr i7_r26_lat_q_7__u1 (.QB (nx8219), .D (nx9340), .CLK (nx2494), .R (
           DecompressedData1[255])) ;
    inv01 i7_r26_lat_q_7__u2 (.Y (DecompressedData1[23]), .A (nx8219)) ;
    buf02 i7_r26_lat_q_7__u3 (.Y (nx5827), .A (nx8219)) ;
    latchr i8_r2_lat_q_7__u1 (.QB (nx8222), .D (nx2692), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_7__u2 (.Y (DecompressedData2[23]), .A (nx8222)) ;
    buf02 i8_r2_lat_q_7__u3 (.Y (nx5829), .A (nx8222)) ;
    latchr i7_r25_lat_q_0__u1 (.QB (nx8225), .D (nx9280), .CLK (nx2708), .R (
           DecompressedData1[255])) ;
    inv01 i7_r25_lat_q_0__u2 (.Y (DecompressedData1[24]), .A (nx8225)) ;
    buf02 i7_r25_lat_q_0__u3 (.Y (nx5833), .A (nx8225)) ;
    latchr i8_r2_lat_q_8__u1 (.QB (nx8228), .D (nx2722), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_8__u2 (.Y (DecompressedData2[24]), .A (nx8228)) ;
    buf02 i8_r2_lat_q_8__u3 (.Y (nx5835), .A (nx8228)) ;
    latchr i7_r25_lat_q_1__u1 (.QB (nx8231), .D (nx9294), .CLK (nx2708), .R (
           DecompressedData1[255])) ;
    inv01 i7_r25_lat_q_1__u2 (.Y (DecompressedData1[25]), .A (nx8231)) ;
    buf02 i7_r25_lat_q_1__u3 (.Y (nx5838), .A (nx8231)) ;
    latchr i8_r2_lat_q_9__u1 (.QB (nx8234), .D (nx2746), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_9__u2 (.Y (DecompressedData2[25]), .A (nx8234)) ;
    buf02 i8_r2_lat_q_9__u3 (.Y (nx5841), .A (nx8234)) ;
    latchr i7_r25_lat_q_2__u1 (.QB (nx8237), .D (nx9304), .CLK (nx2708), .R (
           DecompressedData1[255])) ;
    inv01 i7_r25_lat_q_2__u2 (.Y (DecompressedData1[26]), .A (nx8237)) ;
    buf02 i7_r25_lat_q_2__u3 (.Y (nx5845), .A (nx8237)) ;
    latchr i8_r2_lat_q_10__u1 (.QB (nx8240), .D (nx2770), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_10__u2 (.Y (DecompressedData2[26]), .A (nx8240)) ;
    buf02 i8_r2_lat_q_10__u3 (.Y (nx5847), .A (nx8240)) ;
    latchr i7_r25_lat_q_3__u1 (.QB (nx8243), .D (nx9314), .CLK (nx2708), .R (
           DecompressedData1[255])) ;
    inv01 i7_r25_lat_q_3__u2 (.Y (DecompressedData1[27]), .A (nx8243)) ;
    buf02 i7_r25_lat_q_3__u3 (.Y (nx5850), .A (nx8243)) ;
    latchr i8_r2_lat_q_11__u1 (.QB (nx8246), .D (nx2794), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_11__u2 (.Y (DecompressedData2[27]), .A (nx8246)) ;
    buf02 i8_r2_lat_q_11__u3 (.Y (nx5853), .A (nx8246)) ;
    latchr i7_r25_lat_q_4__u1 (.QB (nx8249), .D (nx9324), .CLK (nx2708), .R (
           DecompressedData1[255])) ;
    inv01 i7_r25_lat_q_4__u2 (.Y (DecompressedData1[28]), .A (nx8249)) ;
    buf02 i7_r25_lat_q_4__u3 (.Y (nx5857), .A (nx8249)) ;
    latchr i8_r2_lat_q_12__u1 (.QB (nx8252), .D (nx2818), .CLK (nx9346), .R (
           DecompressedData1[255])) ;
    inv01 i8_r2_lat_q_12__u2 (.Y (DecompressedData2[28]), .A (nx8252)) ;
    buf02 i8_r2_lat_q_12__u3 (.Y (nx5859), .A (nx8252)) ;
    latchr i7_r24_lat_q_0__u1 (.QB (nx8255), .D (nx9280), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_0__u2 (.Y (DecompressedData1[32]), .A (nx8255)) ;
    buf02 i7_r24_lat_q_0__u3 (.Y (nx5875), .A (nx8255)) ;
    latchr i8_r3_lat_q_0__u1 (.QB (nx8258), .D (nx2914), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_0__u2 (.Y (DecompressedData2[32]), .A (nx8258)) ;
    buf02 i8_r3_lat_q_0__u3 (.Y (nx5877), .A (nx8258)) ;
    latchr i7_r24_lat_q_1__u1 (.QB (nx8261), .D (nx9294), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_1__u2 (.Y (DecompressedData1[33]), .A (nx8261)) ;
    buf02 i7_r24_lat_q_1__u3 (.Y (nx5881), .A (nx8261)) ;
    latchr i8_r3_lat_q_1__u1 (.QB (nx8264), .D (nx2938), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_1__u2 (.Y (DecompressedData2[33]), .A (nx8264)) ;
    buf02 i8_r3_lat_q_1__u3 (.Y (nx5883), .A (nx8264)) ;
    latchr i7_r24_lat_q_2__u1 (.QB (nx8267), .D (nx9304), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_2__u2 (.Y (DecompressedData1[34]), .A (nx8267)) ;
    buf02 i7_r24_lat_q_2__u3 (.Y (nx5886), .A (nx8267)) ;
    latchr i8_r3_lat_q_2__u1 (.QB (nx8270), .D (nx2962), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_2__u2 (.Y (DecompressedData2[34]), .A (nx8270)) ;
    buf02 i8_r3_lat_q_2__u3 (.Y (nx5889), .A (nx8270)) ;
    latchr i7_r24_lat_q_3__u1 (.QB (nx8273), .D (nx9314), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_3__u2 (.Y (DecompressedData1[35]), .A (nx8273)) ;
    buf02 i7_r24_lat_q_3__u3 (.Y (nx5893), .A (nx8273)) ;
    latchr i8_r3_lat_q_3__u1 (.QB (nx8276), .D (nx2986), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_3__u2 (.Y (DecompressedData2[35]), .A (nx8276)) ;
    buf02 i8_r3_lat_q_3__u3 (.Y (nx5895), .A (nx8276)) ;
    latchr i7_r24_lat_q_4__u1 (.QB (nx8279), .D (nx9324), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_4__u2 (.Y (DecompressedData1[36]), .A (nx8279)) ;
    buf02 i7_r24_lat_q_4__u3 (.Y (nx5898), .A (nx8279)) ;
    latchr i8_r3_lat_q_4__u1 (.QB (nx8282), .D (nx3010), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_4__u2 (.Y (DecompressedData2[36]), .A (nx8282)) ;
    buf02 i8_r3_lat_q_4__u3 (.Y (nx5901), .A (nx8282)) ;
    latchr i7_r24_lat_q_5__u1 (.QB (nx8285), .D (nx9332), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_5__u2 (.Y (DecompressedData1[37]), .A (nx8285)) ;
    buf02 i7_r24_lat_q_5__u3 (.Y (nx5905), .A (nx8285)) ;
    latchr i8_r3_lat_q_5__u1 (.QB (nx8288), .D (nx3034), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_5__u2 (.Y (DecompressedData2[37]), .A (nx8288)) ;
    buf02 i8_r3_lat_q_5__u3 (.Y (nx5907), .A (nx8288)) ;
    latchr i7_r24_lat_q_6__u1 (.QB (nx8291), .D (nx9336), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_6__u2 (.Y (DecompressedData1[38]), .A (nx8291)) ;
    buf02 i7_r24_lat_q_6__u3 (.Y (nx5910), .A (nx8291)) ;
    latchr i8_r3_lat_q_6__u1 (.QB (nx8294), .D (nx3058), .CLK (nx9348), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_6__u2 (.Y (DecompressedData2[38]), .A (nx8294)) ;
    buf02 i8_r3_lat_q_6__u3 (.Y (nx5913), .A (nx8294)) ;
    latchr i7_r24_lat_q_7__u1 (.QB (nx8297), .D (nx9340), .CLK (nx2888), .R (
           DecompressedData1[255])) ;
    inv01 i7_r24_lat_q_7__u2 (.Y (DecompressedData1[39]), .A (nx8297)) ;
    buf02 i7_r24_lat_q_7__u3 (.Y (nx5917), .A (nx8297)) ;
    latchr i8_r3_lat_q_7__u1 (.QB (nx8300), .D (nx3082), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_7__u2 (.Y (DecompressedData2[39]), .A (nx8300)) ;
    buf02 i8_r3_lat_q_7__u3 (.Y (nx5919), .A (nx8300)) ;
    latchr i7_r23_lat_q_0__u1 (.QB (nx8303), .D (nx9280), .CLK (nx3098), .R (
           DecompressedData1[255])) ;
    inv01 i7_r23_lat_q_0__u2 (.Y (DecompressedData1[40]), .A (nx8303)) ;
    buf02 i7_r23_lat_q_0__u3 (.Y (nx5922), .A (nx8303)) ;
    latchr i8_r3_lat_q_8__u1 (.QB (nx8306), .D (nx3112), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_8__u2 (.Y (DecompressedData2[40]), .A (nx8306)) ;
    buf02 i8_r3_lat_q_8__u3 (.Y (nx5925), .A (nx8306)) ;
    latchr i7_r23_lat_q_1__u1 (.QB (nx8309), .D (nx9294), .CLK (nx3098), .R (
           DecompressedData1[255])) ;
    inv01 i7_r23_lat_q_1__u2 (.Y (DecompressedData1[41]), .A (nx8309)) ;
    buf02 i7_r23_lat_q_1__u3 (.Y (nx5929), .A (nx8309)) ;
    latchr i8_r3_lat_q_9__u1 (.QB (nx8312), .D (nx3136), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_9__u2 (.Y (DecompressedData2[41]), .A (nx8312)) ;
    buf02 i8_r3_lat_q_9__u3 (.Y (nx5931), .A (nx8312)) ;
    latchr i7_r23_lat_q_2__u1 (.QB (nx8315), .D (nx9304), .CLK (nx3098), .R (
           DecompressedData1[255])) ;
    inv01 i7_r23_lat_q_2__u2 (.Y (DecompressedData1[42]), .A (nx8315)) ;
    buf02 i7_r23_lat_q_2__u3 (.Y (nx5934), .A (nx8315)) ;
    latchr i8_r3_lat_q_10__u1 (.QB (nx8318), .D (nx3160), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_10__u2 (.Y (DecompressedData2[42]), .A (nx8318)) ;
    buf02 i8_r3_lat_q_10__u3 (.Y (nx5937), .A (nx8318)) ;
    latchr i7_r23_lat_q_3__u1 (.QB (nx8321), .D (nx9314), .CLK (nx3098), .R (
           DecompressedData1[255])) ;
    inv01 i7_r23_lat_q_3__u2 (.Y (DecompressedData1[43]), .A (nx8321)) ;
    buf02 i7_r23_lat_q_3__u3 (.Y (nx5941), .A (nx8321)) ;
    latchr i8_r3_lat_q_11__u1 (.QB (nx8324), .D (nx3184), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_11__u2 (.Y (DecompressedData2[43]), .A (nx8324)) ;
    buf02 i8_r3_lat_q_11__u3 (.Y (nx5943), .A (nx8324)) ;
    latchr i7_r23_lat_q_4__u1 (.QB (nx8327), .D (nx9324), .CLK (nx3098), .R (
           DecompressedData1[255])) ;
    inv01 i7_r23_lat_q_4__u2 (.Y (DecompressedData1[44]), .A (nx8327)) ;
    buf02 i7_r23_lat_q_4__u3 (.Y (nx5946), .A (nx8327)) ;
    latchr i8_r3_lat_q_12__u1 (.QB (nx8330), .D (nx3208), .CLK (nx9350), .R (
           DecompressedData1[255])) ;
    inv01 i8_r3_lat_q_12__u2 (.Y (DecompressedData2[44]), .A (nx8330)) ;
    buf02 i8_r3_lat_q_12__u3 (.Y (nx5949), .A (nx8330)) ;
    latchr i7_r22_lat_q_0__u1 (.QB (nx8333), .D (nx9280), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_0__u2 (.Y (DecompressedData1[48]), .A (nx8333)) ;
    buf02 i7_r22_lat_q_0__u3 (.Y (nx5965), .A (nx8333)) ;
    latchr i8_r4_lat_q_0__u1 (.QB (nx8336), .D (nx3302), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_0__u2 (.Y (DecompressedData2[48]), .A (nx8336)) ;
    buf02 i8_r4_lat_q_0__u3 (.Y (nx5967), .A (nx8336)) ;
    latchr i7_r22_lat_q_1__u1 (.QB (nx8339), .D (nx9294), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_1__u2 (.Y (DecompressedData1[49]), .A (nx8339)) ;
    buf02 i7_r22_lat_q_1__u3 (.Y (nx5970), .A (nx8339)) ;
    latchr i8_r4_lat_q_1__u1 (.QB (nx8342), .D (nx3326), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_1__u2 (.Y (DecompressedData2[49]), .A (nx8342)) ;
    buf02 i8_r4_lat_q_1__u3 (.Y (nx5973), .A (nx8342)) ;
    latchr i7_r22_lat_q_2__u1 (.QB (nx8345), .D (nx9304), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_2__u2 (.Y (DecompressedData1[50]), .A (nx8345)) ;
    buf02 i7_r22_lat_q_2__u3 (.Y (nx5977), .A (nx8345)) ;
    latchr i8_r4_lat_q_2__u1 (.QB (nx8348), .D (nx3350), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_2__u2 (.Y (DecompressedData2[50]), .A (nx8348)) ;
    buf02 i8_r4_lat_q_2__u3 (.Y (nx5979), .A (nx8348)) ;
    latchr i7_r22_lat_q_3__u1 (.QB (nx8351), .D (nx9314), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_3__u2 (.Y (DecompressedData1[51]), .A (nx8351)) ;
    buf02 i7_r22_lat_q_3__u3 (.Y (nx5982), .A (nx8351)) ;
    latchr i8_r4_lat_q_3__u1 (.QB (nx8354), .D (nx3374), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_3__u2 (.Y (DecompressedData2[51]), .A (nx8354)) ;
    buf02 i8_r4_lat_q_3__u3 (.Y (nx5985), .A (nx8354)) ;
    latchr i7_r22_lat_q_4__u1 (.QB (nx8357), .D (nx9324), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_4__u2 (.Y (DecompressedData1[52]), .A (nx8357)) ;
    buf02 i7_r22_lat_q_4__u3 (.Y (nx5989), .A (nx8357)) ;
    latchr i8_r4_lat_q_4__u1 (.QB (nx8360), .D (nx3398), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_4__u2 (.Y (DecompressedData2[52]), .A (nx8360)) ;
    buf02 i8_r4_lat_q_4__u3 (.Y (nx5991), .A (nx8360)) ;
    latchr i7_r22_lat_q_5__u1 (.QB (nx8363), .D (nx9332), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_5__u2 (.Y (DecompressedData1[53]), .A (nx8363)) ;
    buf02 i7_r22_lat_q_5__u3 (.Y (nx5994), .A (nx8363)) ;
    latchr i8_r4_lat_q_5__u1 (.QB (nx8366), .D (nx3422), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_5__u2 (.Y (DecompressedData2[53]), .A (nx8366)) ;
    buf02 i8_r4_lat_q_5__u3 (.Y (nx5997), .A (nx8366)) ;
    latchr i7_r22_lat_q_6__u1 (.QB (nx8369), .D (nx9336), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_6__u2 (.Y (DecompressedData1[54]), .A (nx8369)) ;
    buf02 i7_r22_lat_q_6__u3 (.Y (nx6001), .A (nx8369)) ;
    latchr i8_r4_lat_q_6__u1 (.QB (nx8372), .D (nx3446), .CLK (nx9352), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_6__u2 (.Y (DecompressedData2[54]), .A (nx8372)) ;
    buf02 i8_r4_lat_q_6__u3 (.Y (nx6003), .A (nx8372)) ;
    latchr i7_r22_lat_q_7__u1 (.QB (nx8375), .D (nx9340), .CLK (nx3272), .R (
           DecompressedData1[255])) ;
    inv01 i7_r22_lat_q_7__u2 (.Y (DecompressedData1[55]), .A (nx8375)) ;
    buf02 i7_r22_lat_q_7__u3 (.Y (nx6007), .A (nx8375)) ;
    latchr i8_r4_lat_q_7__u1 (.QB (nx8378), .D (nx3470), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_7__u2 (.Y (DecompressedData2[55]), .A (nx8378)) ;
    buf02 i8_r4_lat_q_7__u3 (.Y (nx6009), .A (nx8378)) ;
    latchr i7_r21_lat_q_0__u1 (.QB (nx8381), .D (nx9282), .CLK (nx3486), .R (
           DecompressedData1[255])) ;
    inv01 i7_r21_lat_q_0__u2 (.Y (DecompressedData1[56]), .A (nx8381)) ;
    buf02 i7_r21_lat_q_0__u3 (.Y (nx6013), .A (nx8381)) ;
    latchr i8_r4_lat_q_8__u1 (.QB (nx8384), .D (nx3500), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_8__u2 (.Y (DecompressedData2[56]), .A (nx8384)) ;
    buf02 i8_r4_lat_q_8__u3 (.Y (nx6015), .A (nx8384)) ;
    latchr i7_r21_lat_q_1__u1 (.QB (nx8387), .D (nx9296), .CLK (nx3486), .R (
           DecompressedData1[255])) ;
    inv01 i7_r21_lat_q_1__u2 (.Y (DecompressedData1[57]), .A (nx8387)) ;
    buf02 i7_r21_lat_q_1__u3 (.Y (nx6018), .A (nx8387)) ;
    latchr i8_r4_lat_q_9__u1 (.QB (nx8390), .D (nx3524), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_9__u2 (.Y (DecompressedData2[57]), .A (nx8390)) ;
    buf02 i8_r4_lat_q_9__u3 (.Y (nx6021), .A (nx8390)) ;
    latchr i7_r21_lat_q_2__u1 (.QB (nx8393), .D (nx9306), .CLK (nx3486), .R (
           DecompressedData1[255])) ;
    inv01 i7_r21_lat_q_2__u2 (.Y (DecompressedData1[58]), .A (nx8393)) ;
    buf02 i7_r21_lat_q_2__u3 (.Y (nx6025), .A (nx8393)) ;
    latchr i8_r4_lat_q_10__u1 (.QB (nx8396), .D (nx3548), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_10__u2 (.Y (DecompressedData2[58]), .A (nx8396)) ;
    buf02 i8_r4_lat_q_10__u3 (.Y (nx6027), .A (nx8396)) ;
    latchr i7_r21_lat_q_3__u1 (.QB (nx8399), .D (nx9316), .CLK (nx3486), .R (
           DecompressedData1[255])) ;
    inv01 i7_r21_lat_q_3__u2 (.Y (DecompressedData1[59]), .A (nx8399)) ;
    buf02 i7_r21_lat_q_3__u3 (.Y (nx6031), .A (nx8399)) ;
    latchr i8_r4_lat_q_11__u1 (.QB (nx8402), .D (nx3572), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_11__u2 (.Y (DecompressedData2[59]), .A (nx8402)) ;
    buf02 i8_r4_lat_q_11__u3 (.Y (nx6033), .A (nx8402)) ;
    latchr i7_r21_lat_q_4__u1 (.QB (nx8405), .D (nx9326), .CLK (nx3486), .R (
           DecompressedData1[255])) ;
    inv01 i7_r21_lat_q_4__u2 (.Y (DecompressedData1[60]), .A (nx8405)) ;
    buf02 i7_r21_lat_q_4__u3 (.Y (nx6037), .A (nx8405)) ;
    latchr i8_r4_lat_q_12__u1 (.QB (nx8408), .D (nx3596), .CLK (nx9354), .R (
           DecompressedData1[255])) ;
    inv01 i8_r4_lat_q_12__u2 (.Y (DecompressedData2[60]), .A (nx8408)) ;
    buf02 i8_r4_lat_q_12__u3 (.Y (nx6039), .A (nx8408)) ;
    latchr i7_r20_lat_q_0__u1 (.QB (nx8411), .D (nx9282), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_0__u2 (.Y (DecompressedData1[64]), .A (nx8411)) ;
    buf02 i7_r20_lat_q_0__u3 (.Y (nx6055), .A (nx8411)) ;
    latchr i8_r5_lat_q_0__u1 (.QB (nx8414), .D (nx3702), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_0__u2 (.Y (DecompressedData2[64]), .A (nx8414)) ;
    buf02 i8_r5_lat_q_0__u3 (.Y (nx6057), .A (nx8414)) ;
    latchr i7_r20_lat_q_1__u1 (.QB (nx8417), .D (nx9296), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_1__u2 (.Y (DecompressedData1[65]), .A (nx8417)) ;
    buf02 i7_r20_lat_q_1__u3 (.Y (nx6061), .A (nx8417)) ;
    latchr i8_r5_lat_q_1__u1 (.QB (nx8420), .D (nx3726), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_1__u2 (.Y (DecompressedData2[65]), .A (nx8420)) ;
    buf02 i8_r5_lat_q_1__u3 (.Y (nx6063), .A (nx8420)) ;
    latchr i7_r20_lat_q_2__u1 (.QB (nx8423), .D (nx9306), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_2__u2 (.Y (DecompressedData1[66]), .A (nx8423)) ;
    buf02 i7_r20_lat_q_2__u3 (.Y (nx6066), .A (nx8423)) ;
    latchr i8_r5_lat_q_2__u1 (.QB (nx8426), .D (nx3750), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_2__u2 (.Y (DecompressedData2[66]), .A (nx8426)) ;
    buf02 i8_r5_lat_q_2__u3 (.Y (nx6069), .A (nx8426)) ;
    latchr i7_r20_lat_q_3__u1 (.QB (nx8429), .D (nx9316), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_3__u2 (.Y (DecompressedData1[67]), .A (nx8429)) ;
    buf02 i7_r20_lat_q_3__u3 (.Y (nx6073), .A (nx8429)) ;
    latchr i8_r5_lat_q_3__u1 (.QB (nx8432), .D (nx3774), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_3__u2 (.Y (DecompressedData2[67]), .A (nx8432)) ;
    buf02 i8_r5_lat_q_3__u3 (.Y (nx6075), .A (nx8432)) ;
    latchr i7_r20_lat_q_4__u1 (.QB (nx8435), .D (nx9326), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_4__u2 (.Y (DecompressedData1[68]), .A (nx8435)) ;
    buf02 i7_r20_lat_q_4__u3 (.Y (nx6078), .A (nx8435)) ;
    latchr i8_r5_lat_q_4__u1 (.QB (nx8438), .D (nx3798), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_4__u2 (.Y (DecompressedData2[68]), .A (nx8438)) ;
    buf02 i8_r5_lat_q_4__u3 (.Y (nx6081), .A (nx8438)) ;
    latchr i7_r20_lat_q_5__u1 (.QB (nx8441), .D (nx9332), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_5__u2 (.Y (DecompressedData1[69]), .A (nx8441)) ;
    buf02 i7_r20_lat_q_5__u3 (.Y (nx6085), .A (nx8441)) ;
    latchr i8_r5_lat_q_5__u1 (.QB (nx8444), .D (nx3822), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_5__u2 (.Y (DecompressedData2[69]), .A (nx8444)) ;
    buf02 i8_r5_lat_q_5__u3 (.Y (nx6087), .A (nx8444)) ;
    latchr i7_r20_lat_q_6__u1 (.QB (nx8447), .D (nx9336), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_6__u2 (.Y (DecompressedData1[70]), .A (nx8447)) ;
    buf02 i7_r20_lat_q_6__u3 (.Y (nx6090), .A (nx8447)) ;
    latchr i8_r5_lat_q_6__u1 (.QB (nx8450), .D (nx3846), .CLK (nx9356), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_6__u2 (.Y (DecompressedData2[70]), .A (nx8450)) ;
    buf02 i8_r5_lat_q_6__u3 (.Y (nx6093), .A (nx8450)) ;
    latchr i7_r20_lat_q_7__u1 (.QB (nx8453), .D (nx9340), .CLK (nx3668), .R (
           DecompressedData1[255])) ;
    inv01 i7_r20_lat_q_7__u2 (.Y (DecompressedData1[71]), .A (nx8453)) ;
    buf02 i7_r20_lat_q_7__u3 (.Y (nx6097), .A (nx8453)) ;
    latchr i8_r5_lat_q_7__u1 (.QB (nx8456), .D (nx3870), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_7__u2 (.Y (DecompressedData2[71]), .A (nx8456)) ;
    buf02 i8_r5_lat_q_7__u3 (.Y (nx6099), .A (nx8456)) ;
    latchr i7_r19_lat_q_0__u1 (.QB (nx8459), .D (nx9282), .CLK (nx3886), .R (
           DecompressedData1[255])) ;
    inv01 i7_r19_lat_q_0__u2 (.Y (DecompressedData1[72]), .A (nx8459)) ;
    buf02 i7_r19_lat_q_0__u3 (.Y (nx6102), .A (nx8459)) ;
    latchr i8_r5_lat_q_8__u1 (.QB (nx8462), .D (nx3900), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_8__u2 (.Y (DecompressedData2[72]), .A (nx8462)) ;
    buf02 i8_r5_lat_q_8__u3 (.Y (nx6105), .A (nx8462)) ;
    latchr i7_r19_lat_q_1__u1 (.QB (nx8465), .D (nx9296), .CLK (nx3886), .R (
           DecompressedData1[255])) ;
    inv01 i7_r19_lat_q_1__u2 (.Y (DecompressedData1[73]), .A (nx8465)) ;
    buf02 i7_r19_lat_q_1__u3 (.Y (nx6109), .A (nx8465)) ;
    latchr i8_r5_lat_q_9__u1 (.QB (nx8468), .D (nx3924), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_9__u2 (.Y (DecompressedData2[73]), .A (nx8468)) ;
    buf02 i8_r5_lat_q_9__u3 (.Y (nx6111), .A (nx8468)) ;
    latchr i7_r19_lat_q_2__u1 (.QB (nx8471), .D (nx9306), .CLK (nx3886), .R (
           DecompressedData1[255])) ;
    inv01 i7_r19_lat_q_2__u2 (.Y (DecompressedData1[74]), .A (nx8471)) ;
    buf02 i7_r19_lat_q_2__u3 (.Y (nx6114), .A (nx8471)) ;
    latchr i8_r5_lat_q_10__u1 (.QB (nx8474), .D (nx3948), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_10__u2 (.Y (DecompressedData2[74]), .A (nx8474)) ;
    buf02 i8_r5_lat_q_10__u3 (.Y (nx6117), .A (nx8474)) ;
    latchr i7_r19_lat_q_3__u1 (.QB (nx8477), .D (nx9316), .CLK (nx3886), .R (
           DecompressedData1[255])) ;
    inv01 i7_r19_lat_q_3__u2 (.Y (DecompressedData1[75]), .A (nx8477)) ;
    buf02 i7_r19_lat_q_3__u3 (.Y (nx6121), .A (nx8477)) ;
    latchr i8_r5_lat_q_11__u1 (.QB (nx8480), .D (nx3972), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_11__u2 (.Y (DecompressedData2[75]), .A (nx8480)) ;
    buf02 i8_r5_lat_q_11__u3 (.Y (nx6123), .A (nx8480)) ;
    latchr i7_r19_lat_q_4__u1 (.QB (nx8483), .D (nx9326), .CLK (nx3886), .R (
           DecompressedData1[255])) ;
    inv01 i7_r19_lat_q_4__u2 (.Y (DecompressedData1[76]), .A (nx8483)) ;
    buf02 i7_r19_lat_q_4__u3 (.Y (nx6126), .A (nx8483)) ;
    latchr i8_r5_lat_q_12__u1 (.QB (nx8486), .D (nx3996), .CLK (nx9358), .R (
           DecompressedData1[255])) ;
    inv01 i8_r5_lat_q_12__u2 (.Y (DecompressedData2[76]), .A (nx8486)) ;
    buf02 i8_r5_lat_q_12__u3 (.Y (nx6129), .A (nx8486)) ;
    latchr i7_r18_lat_q_0__u1 (.QB (nx8489), .D (nx9282), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_0__u2 (.Y (DecompressedData1[80]), .A (nx8489)) ;
    buf02 i7_r18_lat_q_0__u3 (.Y (nx6145), .A (nx8489)) ;
    latchr i8_r6_lat_q_0__u1 (.QB (nx8492), .D (nx4086), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_0__u2 (.Y (DecompressedData2[80]), .A (nx8492)) ;
    buf02 i8_r6_lat_q_0__u3 (.Y (nx6147), .A (nx8492)) ;
    latchr i7_r18_lat_q_1__u1 (.QB (nx8495), .D (nx9296), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_1__u2 (.Y (DecompressedData1[81]), .A (nx8495)) ;
    buf02 i7_r18_lat_q_1__u3 (.Y (nx6150), .A (nx8495)) ;
    latchr i8_r6_lat_q_1__u1 (.QB (nx8498), .D (nx4110), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_1__u2 (.Y (DecompressedData2[81]), .A (nx8498)) ;
    buf02 i8_r6_lat_q_1__u3 (.Y (nx6153), .A (nx8498)) ;
    latchr i7_r18_lat_q_2__u1 (.QB (nx8501), .D (nx9306), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_2__u2 (.Y (DecompressedData1[82]), .A (nx8501)) ;
    buf02 i7_r18_lat_q_2__u3 (.Y (nx6157), .A (nx8501)) ;
    latchr i8_r6_lat_q_2__u1 (.QB (nx8504), .D (nx4134), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_2__u2 (.Y (DecompressedData2[82]), .A (nx8504)) ;
    buf02 i8_r6_lat_q_2__u3 (.Y (nx6159), .A (nx8504)) ;
    latchr i7_r18_lat_q_3__u1 (.QB (nx8507), .D (nx9316), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_3__u2 (.Y (DecompressedData1[83]), .A (nx8507)) ;
    buf02 i7_r18_lat_q_3__u3 (.Y (nx6162), .A (nx8507)) ;
    latchr i8_r6_lat_q_3__u1 (.QB (nx8510), .D (nx4158), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_3__u2 (.Y (DecompressedData2[83]), .A (nx8510)) ;
    buf02 i8_r6_lat_q_3__u3 (.Y (nx6165), .A (nx8510)) ;
    latchr i7_r18_lat_q_4__u1 (.QB (nx8513), .D (nx9326), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_4__u2 (.Y (DecompressedData1[84]), .A (nx8513)) ;
    buf02 i7_r18_lat_q_4__u3 (.Y (nx6169), .A (nx8513)) ;
    latchr i8_r6_lat_q_4__u1 (.QB (nx8516), .D (nx4182), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_4__u2 (.Y (DecompressedData2[84]), .A (nx8516)) ;
    buf02 i8_r6_lat_q_4__u3 (.Y (nx6171), .A (nx8516)) ;
    latchr i7_r18_lat_q_5__u1 (.QB (nx8519), .D (nx9332), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_5__u2 (.Y (DecompressedData1[85]), .A (nx8519)) ;
    buf02 i7_r18_lat_q_5__u3 (.Y (nx6174), .A (nx8519)) ;
    latchr i8_r6_lat_q_5__u1 (.QB (nx8522), .D (nx4206), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_5__u2 (.Y (DecompressedData2[85]), .A (nx8522)) ;
    buf02 i8_r6_lat_q_5__u3 (.Y (nx6177), .A (nx8522)) ;
    latchr i7_r18_lat_q_6__u1 (.QB (nx8525), .D (nx9336), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_6__u2 (.Y (DecompressedData1[86]), .A (nx8525)) ;
    buf02 i7_r18_lat_q_6__u3 (.Y (nx6181), .A (nx8525)) ;
    latchr i8_r6_lat_q_6__u1 (.QB (nx8528), .D (nx4230), .CLK (nx9360), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_6__u2 (.Y (DecompressedData2[86]), .A (nx8528)) ;
    buf02 i8_r6_lat_q_6__u3 (.Y (nx6183), .A (nx8528)) ;
    latchr i7_r18_lat_q_7__u1 (.QB (nx8531), .D (nx9340), .CLK (nx4060), .R (
           DecompressedData1[255])) ;
    inv01 i7_r18_lat_q_7__u2 (.Y (DecompressedData1[87]), .A (nx8531)) ;
    buf02 i7_r18_lat_q_7__u3 (.Y (nx6186), .A (nx8531)) ;
    latchr i8_r6_lat_q_7__u1 (.QB (nx8534), .D (nx4254), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_7__u2 (.Y (DecompressedData2[87]), .A (nx8534)) ;
    buf02 i8_r6_lat_q_7__u3 (.Y (nx6189), .A (nx8534)) ;
    latchr i7_r17_lat_q_0__u1 (.QB (nx8537), .D (nx9282), .CLK (nx4270), .R (
           DecompressedData1[255])) ;
    inv01 i7_r17_lat_q_0__u2 (.Y (DecompressedData1[88]), .A (nx8537)) ;
    buf02 i7_r17_lat_q_0__u3 (.Y (nx6193), .A (nx8537)) ;
    latchr i8_r6_lat_q_8__u1 (.QB (nx8540), .D (nx4284), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_8__u2 (.Y (DecompressedData2[88]), .A (nx8540)) ;
    buf02 i8_r6_lat_q_8__u3 (.Y (nx6195), .A (nx8540)) ;
    latchr i7_r17_lat_q_1__u1 (.QB (nx8543), .D (nx9296), .CLK (nx4270), .R (
           DecompressedData1[255])) ;
    inv01 i7_r17_lat_q_1__u2 (.Y (DecompressedData1[89]), .A (nx8543)) ;
    buf02 i7_r17_lat_q_1__u3 (.Y (nx6198), .A (nx8543)) ;
    latchr i8_r6_lat_q_9__u1 (.QB (nx8546), .D (nx4308), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_9__u2 (.Y (DecompressedData2[89]), .A (nx8546)) ;
    buf02 i8_r6_lat_q_9__u3 (.Y (nx6201), .A (nx8546)) ;
    latchr i7_r17_lat_q_2__u1 (.QB (nx8549), .D (nx9306), .CLK (nx4270), .R (
           DecompressedData1[255])) ;
    inv01 i7_r17_lat_q_2__u2 (.Y (DecompressedData1[90]), .A (nx8549)) ;
    buf02 i7_r17_lat_q_2__u3 (.Y (nx6205), .A (nx8549)) ;
    latchr i8_r6_lat_q_10__u1 (.QB (nx8552), .D (nx4332), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_10__u2 (.Y (DecompressedData2[90]), .A (nx8552)) ;
    buf02 i8_r6_lat_q_10__u3 (.Y (nx6207), .A (nx8552)) ;
    latchr i7_r17_lat_q_3__u1 (.QB (nx8555), .D (nx9316), .CLK (nx4270), .R (
           DecompressedData1[255])) ;
    inv01 i7_r17_lat_q_3__u2 (.Y (DecompressedData1[91]), .A (nx8555)) ;
    buf02 i7_r17_lat_q_3__u3 (.Y (nx6210), .A (nx8555)) ;
    latchr i8_r6_lat_q_11__u1 (.QB (nx8558), .D (nx4356), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_11__u2 (.Y (DecompressedData2[91]), .A (nx8558)) ;
    buf02 i8_r6_lat_q_11__u3 (.Y (nx6213), .A (nx8558)) ;
    latchr i7_r17_lat_q_4__u1 (.QB (nx8561), .D (nx9326), .CLK (nx4270), .R (
           DecompressedData1[255])) ;
    inv01 i7_r17_lat_q_4__u2 (.Y (DecompressedData1[92]), .A (nx8561)) ;
    buf02 i7_r17_lat_q_4__u3 (.Y (nx6217), .A (nx8561)) ;
    latchr i8_r6_lat_q_12__u1 (.QB (nx8564), .D (nx4380), .CLK (nx9362), .R (
           DecompressedData1[255])) ;
    inv01 i8_r6_lat_q_12__u2 (.Y (DecompressedData2[92]), .A (nx8564)) ;
    buf02 i8_r6_lat_q_12__u3 (.Y (nx6219), .A (nx8564)) ;
    latchr i7_r16_lat_q_0__u1 (.QB (nx8567), .D (nx9282), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_0__u2 (.Y (DecompressedData1[96]), .A (nx8567)) ;
    buf02 i7_r16_lat_q_0__u3 (.Y (nx6235), .A (nx8567)) ;
    latchr i8_r7_lat_q_0__u1 (.QB (nx8570), .D (nx4480), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_0__u2 (.Y (DecompressedData2[96]), .A (nx8570)) ;
    buf02 i8_r7_lat_q_0__u3 (.Y (nx6237), .A (nx8570)) ;
    latchr i7_r16_lat_q_1__u1 (.QB (nx8573), .D (nx9296), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_1__u2 (.Y (DecompressedData1[97]), .A (nx8573)) ;
    buf02 i7_r16_lat_q_1__u3 (.Y (nx6240), .A (nx8573)) ;
    latchr i8_r7_lat_q_1__u1 (.QB (nx8576), .D (nx4504), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_1__u2 (.Y (DecompressedData2[97]), .A (nx8576)) ;
    buf02 i8_r7_lat_q_1__u3 (.Y (nx6243), .A (nx8576)) ;
    latchr i7_r16_lat_q_2__u1 (.QB (nx8579), .D (nx9306), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_2__u2 (.Y (DecompressedData1[98]), .A (nx8579)) ;
    buf02 i7_r16_lat_q_2__u3 (.Y (nx6247), .A (nx8579)) ;
    latchr i8_r7_lat_q_2__u1 (.QB (nx8582), .D (nx4528), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_2__u2 (.Y (DecompressedData2[98]), .A (nx8582)) ;
    buf02 i8_r7_lat_q_2__u3 (.Y (nx6249), .A (nx8582)) ;
    latchr i7_r16_lat_q_3__u1 (.QB (nx8585), .D (nx9316), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_3__u2 (.Y (DecompressedData1[99]), .A (nx8585)) ;
    buf02 i7_r16_lat_q_3__u3 (.Y (nx6252), .A (nx8585)) ;
    latchr i8_r7_lat_q_3__u1 (.QB (nx8588), .D (nx4552), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_3__u2 (.Y (DecompressedData2[99]), .A (nx8588)) ;
    buf02 i8_r7_lat_q_3__u3 (.Y (nx6255), .A (nx8588)) ;
    latchr i7_r16_lat_q_4__u1 (.QB (nx8591), .D (nx9326), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_4__u2 (.Y (DecompressedData1[100]), .A (nx8591)) ;
    buf02 i7_r16_lat_q_4__u3 (.Y (nx6259), .A (nx8591)) ;
    latchr i8_r7_lat_q_4__u1 (.QB (nx8594), .D (nx4576), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_4__u2 (.Y (DecompressedData2[100]), .A (nx8594)) ;
    buf02 i8_r7_lat_q_4__u3 (.Y (nx6261), .A (nx8594)) ;
    latchr i7_r16_lat_q_5__u1 (.QB (nx8597), .D (nx9332), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_5__u2 (.Y (DecompressedData1[101]), .A (nx8597)) ;
    buf02 i7_r16_lat_q_5__u3 (.Y (nx6264), .A (nx8597)) ;
    latchr i8_r7_lat_q_5__u1 (.QB (nx8600), .D (nx4600), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_5__u2 (.Y (DecompressedData2[101]), .A (nx8600)) ;
    buf02 i8_r7_lat_q_5__u3 (.Y (nx6267), .A (nx8600)) ;
    latchr i7_r16_lat_q_6__u1 (.QB (nx8603), .D (nx9336), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_6__u2 (.Y (DecompressedData1[102]), .A (nx8603)) ;
    buf02 i7_r16_lat_q_6__u3 (.Y (nx6271), .A (nx8603)) ;
    latchr i8_r7_lat_q_6__u1 (.QB (nx8606), .D (nx4624), .CLK (nx9364), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_6__u2 (.Y (DecompressedData2[102]), .A (nx8606)) ;
    buf02 i8_r7_lat_q_6__u3 (.Y (nx6273), .A (nx8606)) ;
    latchr i7_r16_lat_q_7__u1 (.QB (nx8609), .D (nx9340), .CLK (nx4454), .R (
           DecompressedData1[255])) ;
    inv01 i7_r16_lat_q_7__u2 (.Y (DecompressedData1[103]), .A (nx8609)) ;
    buf02 i7_r16_lat_q_7__u3 (.Y (nx6276), .A (nx8609)) ;
    latchr i8_r7_lat_q_7__u1 (.QB (nx8612), .D (nx4648), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_7__u2 (.Y (DecompressedData2[103]), .A (nx8612)) ;
    buf02 i8_r7_lat_q_7__u3 (.Y (nx6279), .A (nx8612)) ;
    latchr i7_r15_lat_q_0__u1 (.QB (nx8615), .D (nx9282), .CLK (nx4664), .R (
           DecompressedData1[255])) ;
    inv01 i7_r15_lat_q_0__u2 (.Y (DecompressedData1[104]), .A (nx8615)) ;
    buf02 i7_r15_lat_q_0__u3 (.Y (nx6283), .A (nx8615)) ;
    latchr i8_r7_lat_q_8__u1 (.QB (nx8618), .D (nx4678), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_8__u2 (.Y (DecompressedData2[104]), .A (nx8618)) ;
    buf02 i8_r7_lat_q_8__u3 (.Y (nx6285), .A (nx8618)) ;
    latchr i7_r15_lat_q_1__u1 (.QB (nx8621), .D (nx9296), .CLK (nx4664), .R (
           DecompressedData1[255])) ;
    inv01 i7_r15_lat_q_1__u2 (.Y (DecompressedData1[105]), .A (nx8621)) ;
    buf02 i7_r15_lat_q_1__u3 (.Y (nx6288), .A (nx8621)) ;
    latchr i8_r7_lat_q_9__u1 (.QB (nx8624), .D (nx4702), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_9__u2 (.Y (DecompressedData2[105]), .A (nx8624)) ;
    buf02 i8_r7_lat_q_9__u3 (.Y (nx6291), .A (nx8624)) ;
    latchr i7_r15_lat_q_2__u1 (.QB (nx8627), .D (nx9306), .CLK (nx4664), .R (
           DecompressedData1[255])) ;
    inv01 i7_r15_lat_q_2__u2 (.Y (DecompressedData1[106]), .A (nx8627)) ;
    buf02 i7_r15_lat_q_2__u3 (.Y (nx6295), .A (nx8627)) ;
    latchr i8_r7_lat_q_10__u1 (.QB (nx8630), .D (nx4726), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_10__u2 (.Y (DecompressedData2[106]), .A (nx8630)) ;
    buf02 i8_r7_lat_q_10__u3 (.Y (nx6297), .A (nx8630)) ;
    latchr i7_r15_lat_q_3__u1 (.QB (nx8633), .D (nx9316), .CLK (nx4664), .R (
           DecompressedData1[255])) ;
    inv01 i7_r15_lat_q_3__u2 (.Y (DecompressedData1[107]), .A (nx8633)) ;
    buf02 i7_r15_lat_q_3__u3 (.Y (nx6300), .A (nx8633)) ;
    latchr i8_r7_lat_q_11__u1 (.QB (nx8636), .D (nx4750), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_11__u2 (.Y (DecompressedData2[107]), .A (nx8636)) ;
    buf02 i8_r7_lat_q_11__u3 (.Y (nx6303), .A (nx8636)) ;
    latchr i7_r15_lat_q_4__u1 (.QB (nx8639), .D (nx9326), .CLK (nx4664), .R (
           DecompressedData1[255])) ;
    inv01 i7_r15_lat_q_4__u2 (.Y (DecompressedData1[108]), .A (nx8639)) ;
    buf02 i7_r15_lat_q_4__u3 (.Y (nx6307), .A (nx8639)) ;
    latchr i8_r7_lat_q_12__u1 (.QB (nx8642), .D (nx4774), .CLK (nx9366), .R (
           DecompressedData1[255])) ;
    inv01 i8_r7_lat_q_12__u2 (.Y (DecompressedData2[108]), .A (nx8642)) ;
    buf02 i8_r7_lat_q_12__u3 (.Y (nx6309), .A (nx8642)) ;
    latchr i7_r14_lat_q_0__u1 (.QB (nx8645), .D (nx9284), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_0__u2 (.Y (DecompressedData1[112]), .A (nx8645)) ;
    buf02 i7_r14_lat_q_0__u3 (.Y (nx6325), .A (nx8645)) ;
    latchr i8_r8_lat_q_0__u1 (.QB (nx8648), .D (nx4864), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_0__u2 (.Y (DecompressedData2[112]), .A (nx8648)) ;
    buf02 i8_r8_lat_q_0__u3 (.Y (nx6327), .A (nx8648)) ;
    latchr i7_r14_lat_q_1__u1 (.QB (nx8651), .D (nx9298), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_1__u2 (.Y (DecompressedData1[113]), .A (nx8651)) ;
    buf02 i7_r14_lat_q_1__u3 (.Y (nx6331), .A (nx8651)) ;
    latchr i8_r8_lat_q_1__u1 (.QB (nx8654), .D (nx4888), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_1__u2 (.Y (DecompressedData2[113]), .A (nx8654)) ;
    buf02 i8_r8_lat_q_1__u3 (.Y (nx6333), .A (nx8654)) ;
    latchr i7_r14_lat_q_2__u1 (.QB (nx8657), .D (nx9308), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_2__u2 (.Y (DecompressedData1[114]), .A (nx8657)) ;
    buf02 i7_r14_lat_q_2__u3 (.Y (nx6336), .A (nx8657)) ;
    latchr i8_r8_lat_q_2__u1 (.QB (nx8660), .D (nx4912), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_2__u2 (.Y (DecompressedData2[114]), .A (nx8660)) ;
    buf02 i8_r8_lat_q_2__u3 (.Y (nx6339), .A (nx8660)) ;
    latchr i7_r14_lat_q_3__u1 (.QB (nx8663), .D (nx9318), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_3__u2 (.Y (DecompressedData1[115]), .A (nx8663)) ;
    buf02 i7_r14_lat_q_3__u3 (.Y (nx6343), .A (nx8663)) ;
    latchr i8_r8_lat_q_3__u1 (.QB (nx8666), .D (nx4936), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_3__u2 (.Y (DecompressedData2[115]), .A (nx8666)) ;
    buf02 i8_r8_lat_q_3__u3 (.Y (nx6345), .A (nx8666)) ;
    latchr i7_r14_lat_q_4__u1 (.QB (nx8669), .D (nx9328), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_4__u2 (.Y (DecompressedData1[116]), .A (nx8669)) ;
    buf02 i7_r14_lat_q_4__u3 (.Y (nx6348), .A (nx8669)) ;
    latchr i8_r8_lat_q_4__u1 (.QB (nx8672), .D (nx4960), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_4__u2 (.Y (DecompressedData2[116]), .A (nx8672)) ;
    buf02 i8_r8_lat_q_4__u3 (.Y (nx6350), .A (nx8672)) ;
    latchr i7_r14_lat_q_5__u1 (.QB (nx8675), .D (nx9334), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_5__u2 (.Y (DecompressedData1[117]), .A (nx8675)) ;
    buf02 i7_r14_lat_q_5__u3 (.Y (nx6353), .A (nx8675)) ;
    latchr i8_r8_lat_q_5__u1 (.QB (nx8678), .D (nx4984), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_5__u2 (.Y (DecompressedData2[117]), .A (nx8678)) ;
    buf02 i8_r8_lat_q_5__u3 (.Y (nx6355), .A (nx8678)) ;
    latchr i7_r14_lat_q_6__u1 (.QB (nx8681), .D (nx9338), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_6__u2 (.Y (DecompressedData1[118]), .A (nx8681)) ;
    buf02 i7_r14_lat_q_6__u3 (.Y (nx6358), .A (nx8681)) ;
    latchr i8_r8_lat_q_6__u1 (.QB (nx8684), .D (nx5008), .CLK (nx9368), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_6__u2 (.Y (DecompressedData2[118]), .A (nx8684)) ;
    buf02 i8_r8_lat_q_6__u3 (.Y (nx6360), .A (nx8684)) ;
    latchr i7_r14_lat_q_7__u1 (.QB (nx8687), .D (nx9342), .CLK (nx4838), .R (
           DecompressedData1[255])) ;
    inv01 i7_r14_lat_q_7__u2 (.Y (DecompressedData1[119]), .A (nx8687)) ;
    buf02 i7_r14_lat_q_7__u3 (.Y (nx6363), .A (nx8687)) ;
    latchr i8_r8_lat_q_7__u1 (.QB (nx8690), .D (nx5032), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_7__u2 (.Y (DecompressedData2[119]), .A (nx8690)) ;
    buf02 i8_r8_lat_q_7__u3 (.Y (nx6365), .A (nx8690)) ;
    latchr i7_r13_lat_q_0__u1 (.QB (nx8693), .D (nx9284), .CLK (nx5048), .R (
           DecompressedData1[255])) ;
    inv01 i7_r13_lat_q_0__u2 (.Y (DecompressedData1[120]), .A (nx8693)) ;
    buf02 i7_r13_lat_q_0__u3 (.Y (nx6368), .A (nx8693)) ;
    latchr i8_r8_lat_q_8__u1 (.QB (nx8696), .D (nx5062), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_8__u2 (.Y (DecompressedData2[120]), .A (nx8696)) ;
    buf02 i8_r8_lat_q_8__u3 (.Y (nx6370), .A (nx8696)) ;
    latchr i7_r13_lat_q_1__u1 (.QB (nx8699), .D (nx9298), .CLK (nx5048), .R (
           DecompressedData1[255])) ;
    inv01 i7_r13_lat_q_1__u2 (.Y (DecompressedData1[121]), .A (nx8699)) ;
    buf02 i7_r13_lat_q_1__u3 (.Y (nx6373), .A (nx8699)) ;
    latchr i8_r8_lat_q_9__u1 (.QB (nx8702), .D (nx5086), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_9__u2 (.Y (DecompressedData2[121]), .A (nx8702)) ;
    buf02 i8_r8_lat_q_9__u3 (.Y (nx6375), .A (nx8702)) ;
    latchr i7_r13_lat_q_2__u1 (.QB (nx8705), .D (nx9308), .CLK (nx5048), .R (
           DecompressedData1[255])) ;
    inv01 i7_r13_lat_q_2__u2 (.Y (DecompressedData1[122]), .A (nx8705)) ;
    buf02 i7_r13_lat_q_2__u3 (.Y (nx6379), .A (nx8705)) ;
    latchr i8_r8_lat_q_10__u1 (.QB (nx8708), .D (nx5110), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_10__u2 (.Y (DecompressedData2[122]), .A (nx8708)) ;
    buf02 i8_r8_lat_q_10__u3 (.Y (nx6381), .A (nx8708)) ;
    latchr i7_r13_lat_q_3__u1 (.QB (nx8711), .D (nx9318), .CLK (nx5048), .R (
           DecompressedData1[255])) ;
    inv01 i7_r13_lat_q_3__u2 (.Y (DecompressedData1[123]), .A (nx8711)) ;
    buf02 i7_r13_lat_q_3__u3 (.Y (nx6384), .A (nx8711)) ;
    latchr i8_r8_lat_q_11__u1 (.QB (nx8714), .D (nx5134), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_11__u2 (.Y (DecompressedData2[123]), .A (nx8714)) ;
    buf02 i8_r8_lat_q_11__u3 (.Y (nx6387), .A (nx8714)) ;
    latchr i7_r13_lat_q_4__u1 (.QB (nx8717), .D (nx9328), .CLK (nx5048), .R (
           DecompressedData1[255])) ;
    inv01 i7_r13_lat_q_4__u2 (.Y (DecompressedData1[124]), .A (nx8717)) ;
    buf02 i7_r13_lat_q_4__u3 (.Y (nx6391), .A (nx8717)) ;
    latchr i8_r8_lat_q_12__u1 (.QB (nx8720), .D (nx5158), .CLK (nx9370), .R (
           DecompressedData1[255])) ;
    inv01 i8_r8_lat_q_12__u2 (.Y (DecompressedData2[124]), .A (nx8720)) ;
    buf02 i8_r8_lat_q_12__u3 (.Y (nx6393), .A (nx8720)) ;
    latchr i7_r12_lat_q_0__u1 (.QB (nx8723), .D (nx9284), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_0__u2 (.Y (DecompressedData1[128]), .A (nx8723)) ;
    buf02 i7_r12_lat_q_0__u3 (.Y (nx6409), .A (nx8723)) ;
    latchr i8_r9_lat_q_0__u1 (.QB (nx8726), .D (nx5262), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_0__u2 (.Y (DecompressedData2[128]), .A (nx8726)) ;
    buf02 i8_r9_lat_q_0__u3 (.Y (nx6411), .A (nx8726)) ;
    latchr i7_r12_lat_q_1__u1 (.QB (nx8729), .D (nx9298), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_1__u2 (.Y (DecompressedData1[129]), .A (nx8729)) ;
    buf02 i7_r12_lat_q_1__u3 (.Y (nx6415), .A (nx8729)) ;
    latchr i8_r9_lat_q_1__u1 (.QB (nx8732), .D (nx5286), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_1__u2 (.Y (DecompressedData2[129]), .A (nx8732)) ;
    buf02 i8_r9_lat_q_1__u3 (.Y (nx6417), .A (nx8732)) ;
    latchr i7_r12_lat_q_2__u1 (.QB (nx8735), .D (nx9308), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_2__u2 (.Y (DecompressedData1[130]), .A (nx8735)) ;
    buf02 i7_r12_lat_q_2__u3 (.Y (nx6421), .A (nx8735)) ;
    latchr i8_r9_lat_q_2__u1 (.QB (nx8738), .D (nx5310), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_2__u2 (.Y (DecompressedData2[130]), .A (nx8738)) ;
    buf02 i8_r9_lat_q_2__u3 (.Y (nx6423), .A (nx8738)) ;
    latchr i7_r12_lat_q_3__u1 (.QB (nx8741), .D (nx9318), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_3__u2 (.Y (DecompressedData1[131]), .A (nx8741)) ;
    buf02 i7_r12_lat_q_3__u3 (.Y (nx6426), .A (nx8741)) ;
    latchr i8_r9_lat_q_3__u1 (.QB (nx8744), .D (nx5334), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_3__u2 (.Y (DecompressedData2[131]), .A (nx8744)) ;
    buf02 i8_r9_lat_q_3__u3 (.Y (nx6429), .A (nx8744)) ;
    latchr i7_r12_lat_q_4__u1 (.QB (nx8747), .D (nx9328), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_4__u2 (.Y (DecompressedData1[132]), .A (nx8747)) ;
    buf02 i7_r12_lat_q_4__u3 (.Y (nx6433), .A (nx8747)) ;
    latchr i8_r9_lat_q_4__u1 (.QB (nx8750), .D (nx5358), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_4__u2 (.Y (DecompressedData2[132]), .A (nx8750)) ;
    buf02 i8_r9_lat_q_4__u3 (.Y (nx6435), .A (nx8750)) ;
    latchr i7_r12_lat_q_5__u1 (.QB (nx8753), .D (nx9334), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_5__u2 (.Y (DecompressedData1[133]), .A (nx8753)) ;
    buf02 i7_r12_lat_q_5__u3 (.Y (nx6438), .A (nx8753)) ;
    latchr i8_r9_lat_q_5__u1 (.QB (nx8756), .D (nx5382), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_5__u2 (.Y (DecompressedData2[133]), .A (nx8756)) ;
    buf02 i8_r9_lat_q_5__u3 (.Y (nx6441), .A (nx8756)) ;
    latchr i7_r12_lat_q_6__u1 (.QB (nx8759), .D (nx9338), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_6__u2 (.Y (DecompressedData1[134]), .A (nx8759)) ;
    buf02 i7_r12_lat_q_6__u3 (.Y (nx6445), .A (nx8759)) ;
    latchr i8_r9_lat_q_6__u1 (.QB (nx8762), .D (nx5406), .CLK (nx9372), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_6__u2 (.Y (DecompressedData2[134]), .A (nx8762)) ;
    buf02 i8_r9_lat_q_6__u3 (.Y (nx6447), .A (nx8762)) ;
    latchr i7_r12_lat_q_7__u1 (.QB (nx8765), .D (nx9342), .CLK (nx5228), .R (
           DecompressedData1[255])) ;
    inv01 i7_r12_lat_q_7__u2 (.Y (DecompressedData1[135]), .A (nx8765)) ;
    buf02 i7_r12_lat_q_7__u3 (.Y (nx6450), .A (nx8765)) ;
    latchr i8_r9_lat_q_7__u1 (.QB (nx8768), .D (nx5430), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_7__u2 (.Y (DecompressedData2[135]), .A (nx8768)) ;
    buf02 i8_r9_lat_q_7__u3 (.Y (nx6453), .A (nx8768)) ;
    latchr i7_r11_lat_q_0__u1 (.QB (nx8771), .D (nx9284), .CLK (nx5446), .R (
           DecompressedData1[255])) ;
    inv01 i7_r11_lat_q_0__u2 (.Y (DecompressedData1[136]), .A (nx8771)) ;
    buf02 i7_r11_lat_q_0__u3 (.Y (nx6457), .A (nx8771)) ;
    latchr i8_r9_lat_q_8__u1 (.QB (nx8774), .D (nx5460), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_8__u2 (.Y (DecompressedData2[136]), .A (nx8774)) ;
    buf02 i8_r9_lat_q_8__u3 (.Y (nx6459), .A (nx8774)) ;
    latchr i7_r11_lat_q_1__u1 (.QB (nx8777), .D (nx9298), .CLK (nx5446), .R (
           DecompressedData1[255])) ;
    inv01 i7_r11_lat_q_1__u2 (.Y (DecompressedData1[137]), .A (nx8777)) ;
    buf02 i7_r11_lat_q_1__u3 (.Y (nx6462), .A (nx8777)) ;
    latchr i8_r9_lat_q_9__u1 (.QB (nx8780), .D (nx5484), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_9__u2 (.Y (DecompressedData2[137]), .A (nx8780)) ;
    buf02 i8_r9_lat_q_9__u3 (.Y (nx6465), .A (nx8780)) ;
    latchr i7_r11_lat_q_2__u1 (.QB (nx8783), .D (nx9308), .CLK (nx5446), .R (
           DecompressedData1[255])) ;
    inv01 i7_r11_lat_q_2__u2 (.Y (DecompressedData1[138]), .A (nx8783)) ;
    buf02 i7_r11_lat_q_2__u3 (.Y (nx6469), .A (nx8783)) ;
    latchr i8_r9_lat_q_10__u1 (.QB (nx8786), .D (nx5508), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_10__u2 (.Y (DecompressedData2[138]), .A (nx8786)) ;
    buf02 i8_r9_lat_q_10__u3 (.Y (nx6471), .A (nx8786)) ;
    latchr i7_r11_lat_q_3__u1 (.QB (nx8789), .D (nx9318), .CLK (nx5446), .R (
           DecompressedData1[255])) ;
    inv01 i7_r11_lat_q_3__u2 (.Y (DecompressedData1[139]), .A (nx8789)) ;
    buf02 i7_r11_lat_q_3__u3 (.Y (nx6474), .A (nx8789)) ;
    latchr i8_r9_lat_q_11__u1 (.QB (nx8792), .D (nx5532), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_11__u2 (.Y (DecompressedData2[139]), .A (nx8792)) ;
    buf02 i8_r9_lat_q_11__u3 (.Y (nx6477), .A (nx8792)) ;
    latchr i7_r11_lat_q_4__u1 (.QB (nx8795), .D (nx9328), .CLK (nx5446), .R (
           DecompressedData1[255])) ;
    inv01 i7_r11_lat_q_4__u2 (.Y (DecompressedData1[140]), .A (nx8795)) ;
    buf02 i7_r11_lat_q_4__u3 (.Y (nx6481), .A (nx8795)) ;
    latchr i8_r9_lat_q_12__u1 (.QB (nx8798), .D (nx5556), .CLK (nx9374), .R (
           DecompressedData1[255])) ;
    inv01 i8_r9_lat_q_12__u2 (.Y (DecompressedData2[140]), .A (nx8798)) ;
    buf02 i8_r9_lat_q_12__u3 (.Y (nx6483), .A (nx8798)) ;
    latchr i7_r10_lat_q_0__u1 (.QB (nx8801), .D (nx9284), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_0__u2 (.Y (DecompressedData1[144]), .A (nx8801)) ;
    buf02 i7_r10_lat_q_0__u3 (.Y (nx6499), .A (nx8801)) ;
    latchr i8_r10_lat_q_0__u1 (.QB (nx8804), .D (nx5646), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_0__u2 (.Y (DecompressedData2[144]), .A (nx8804)) ;
    buf02 i8_r10_lat_q_0__u3 (.Y (nx6501), .A (nx8804)) ;
    latchr i7_r10_lat_q_1__u1 (.QB (nx8807), .D (nx9298), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_1__u2 (.Y (DecompressedData1[145]), .A (nx8807)) ;
    buf02 i7_r10_lat_q_1__u3 (.Y (nx6505), .A (nx8807)) ;
    latchr i8_r10_lat_q_1__u1 (.QB (nx8810), .D (nx5670), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_1__u2 (.Y (DecompressedData2[145]), .A (nx8810)) ;
    buf02 i8_r10_lat_q_1__u3 (.Y (nx6507), .A (nx8810)) ;
    latchr i7_r10_lat_q_2__u1 (.QB (nx8813), .D (nx9308), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_2__u2 (.Y (DecompressedData1[146]), .A (nx8813)) ;
    buf02 i7_r10_lat_q_2__u3 (.Y (nx6510), .A (nx8813)) ;
    latchr i8_r10_lat_q_2__u1 (.QB (nx8816), .D (nx5694), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_2__u2 (.Y (DecompressedData2[146]), .A (nx8816)) ;
    buf02 i8_r10_lat_q_2__u3 (.Y (nx6513), .A (nx8816)) ;
    latchr i7_r10_lat_q_3__u1 (.QB (nx8819), .D (nx9318), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_3__u2 (.Y (DecompressedData1[147]), .A (nx8819)) ;
    buf02 i7_r10_lat_q_3__u3 (.Y (nx6517), .A (nx8819)) ;
    latchr i8_r10_lat_q_3__u1 (.QB (nx8822), .D (nx5718), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_3__u2 (.Y (DecompressedData2[147]), .A (nx8822)) ;
    buf02 i8_r10_lat_q_3__u3 (.Y (nx6519), .A (nx8822)) ;
    latchr i7_r10_lat_q_4__u1 (.QB (nx8825), .D (nx9328), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_4__u2 (.Y (DecompressedData1[148]), .A (nx8825)) ;
    buf02 i7_r10_lat_q_4__u3 (.Y (nx6522), .A (nx8825)) ;
    latchr i8_r10_lat_q_4__u1 (.QB (nx8828), .D (nx5742), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_4__u2 (.Y (DecompressedData2[148]), .A (nx8828)) ;
    buf02 i8_r10_lat_q_4__u3 (.Y (nx6525), .A (nx8828)) ;
    latchr i7_r10_lat_q_5__u1 (.QB (nx8831), .D (nx9334), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_5__u2 (.Y (DecompressedData1[149]), .A (nx8831)) ;
    buf02 i7_r10_lat_q_5__u3 (.Y (nx6529), .A (nx8831)) ;
    latchr i8_r10_lat_q_5__u1 (.QB (nx8834), .D (nx5766), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_5__u2 (.Y (DecompressedData2[149]), .A (nx8834)) ;
    buf02 i8_r10_lat_q_5__u3 (.Y (nx6531), .A (nx8834)) ;
    latchr i7_r10_lat_q_6__u1 (.QB (nx8837), .D (nx9338), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_6__u2 (.Y (DecompressedData1[150]), .A (nx8837)) ;
    buf02 i7_r10_lat_q_6__u3 (.Y (nx6534), .A (nx8837)) ;
    latchr i8_r10_lat_q_6__u1 (.QB (nx8840), .D (nx5790), .CLK (nx9376), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_6__u2 (.Y (DecompressedData2[150]), .A (nx8840)) ;
    buf02 i8_r10_lat_q_6__u3 (.Y (nx6537), .A (nx8840)) ;
    latchr i7_r10_lat_q_7__u1 (.QB (nx8843), .D (nx9342), .CLK (nx5620), .R (
           DecompressedData1[255])) ;
    inv01 i7_r10_lat_q_7__u2 (.Y (DecompressedData1[151]), .A (nx8843)) ;
    buf02 i7_r10_lat_q_7__u3 (.Y (nx6541), .A (nx8843)) ;
    latchr i8_r10_lat_q_7__u1 (.QB (nx8846), .D (nx5814), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_7__u2 (.Y (DecompressedData2[151]), .A (nx8846)) ;
    buf02 i8_r10_lat_q_7__u3 (.Y (nx6543), .A (nx8846)) ;
    latchr i7_r9_lat_q_0__u1 (.QB (nx8849), .D (nx9284), .CLK (nx5830), .R (
           DecompressedData1[255])) ;
    inv01 i7_r9_lat_q_0__u2 (.Y (DecompressedData1[152]), .A (nx8849)) ;
    buf02 i7_r9_lat_q_0__u3 (.Y (nx6546), .A (nx8849)) ;
    latchr i8_r10_lat_q_8__u1 (.QB (nx8852), .D (nx5844), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_8__u2 (.Y (DecompressedData2[152]), .A (nx8852)) ;
    buf02 i8_r10_lat_q_8__u3 (.Y (nx6549), .A (nx8852)) ;
    latchr i7_r9_lat_q_1__u1 (.QB (nx8855), .D (nx9298), .CLK (nx5830), .R (
           DecompressedData1[255])) ;
    inv01 i7_r9_lat_q_1__u2 (.Y (DecompressedData1[153]), .A (nx8855)) ;
    buf02 i7_r9_lat_q_1__u3 (.Y (nx6553), .A (nx8855)) ;
    latchr i8_r10_lat_q_9__u1 (.QB (nx8858), .D (nx5868), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_9__u2 (.Y (DecompressedData2[153]), .A (nx8858)) ;
    buf02 i8_r10_lat_q_9__u3 (.Y (nx6555), .A (nx8858)) ;
    latchr i7_r9_lat_q_2__u1 (.QB (nx8861), .D (nx9308), .CLK (nx5830), .R (
           DecompressedData1[255])) ;
    inv01 i7_r9_lat_q_2__u2 (.Y (DecompressedData1[154]), .A (nx8861)) ;
    buf02 i7_r9_lat_q_2__u3 (.Y (nx6558), .A (nx8861)) ;
    latchr i8_r10_lat_q_10__u1 (.QB (nx8864), .D (nx5892), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_10__u2 (.Y (DecompressedData2[154]), .A (nx8864)) ;
    buf02 i8_r10_lat_q_10__u3 (.Y (nx6561), .A (nx8864)) ;
    latchr i7_r9_lat_q_3__u1 (.QB (nx8867), .D (nx9318), .CLK (nx5830), .R (
           DecompressedData1[255])) ;
    inv01 i7_r9_lat_q_3__u2 (.Y (DecompressedData1[155]), .A (nx8867)) ;
    buf02 i7_r9_lat_q_3__u3 (.Y (nx6565), .A (nx8867)) ;
    latchr i8_r10_lat_q_11__u1 (.QB (nx8870), .D (nx5916), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_11__u2 (.Y (DecompressedData2[155]), .A (nx8870)) ;
    buf02 i8_r10_lat_q_11__u3 (.Y (nx6567), .A (nx8870)) ;
    latchr i7_r9_lat_q_4__u1 (.QB (nx8873), .D (nx9328), .CLK (nx5830), .R (
           DecompressedData1[255])) ;
    inv01 i7_r9_lat_q_4__u2 (.Y (DecompressedData1[156]), .A (nx8873)) ;
    buf02 i7_r9_lat_q_4__u3 (.Y (nx6570), .A (nx8873)) ;
    latchr i8_r10_lat_q_12__u1 (.QB (nx8876), .D (nx5940), .CLK (nx9378), .R (
           DecompressedData1[255])) ;
    inv01 i8_r10_lat_q_12__u2 (.Y (DecompressedData2[156]), .A (nx8876)) ;
    buf02 i8_r10_lat_q_12__u3 (.Y (nx6573), .A (nx8876)) ;
    latchr i7_r8_lat_q_0__u1 (.QB (nx8879), .D (nx9284), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_0__u2 (.Y (DecompressedData1[160]), .A (nx8879)) ;
    buf02 i7_r8_lat_q_0__u3 (.Y (nx6589), .A (nx8879)) ;
    latchr i8_r11_lat_q_0__u1 (.QB (nx8882), .D (nx6036), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_0__u2 (.Y (DecompressedData2[160]), .A (nx8882)) ;
    buf02 i8_r11_lat_q_0__u3 (.Y (nx6591), .A (nx8882)) ;
    latchr i7_r8_lat_q_1__u1 (.QB (nx8885), .D (nx9298), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_1__u2 (.Y (DecompressedData1[161]), .A (nx8885)) ;
    buf02 i7_r8_lat_q_1__u3 (.Y (nx6594), .A (nx8885)) ;
    latchr i8_r11_lat_q_1__u1 (.QB (nx8888), .D (nx6060), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_1__u2 (.Y (DecompressedData2[161]), .A (nx8888)) ;
    buf02 i8_r11_lat_q_1__u3 (.Y (nx6597), .A (nx8888)) ;
    latchr i7_r8_lat_q_2__u1 (.QB (nx8891), .D (nx9308), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_2__u2 (.Y (DecompressedData1[162]), .A (nx8891)) ;
    buf02 i7_r8_lat_q_2__u3 (.Y (nx6601), .A (nx8891)) ;
    latchr i8_r11_lat_q_2__u1 (.QB (nx8894), .D (nx6084), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_2__u2 (.Y (DecompressedData2[162]), .A (nx8894)) ;
    buf02 i8_r11_lat_q_2__u3 (.Y (nx6603), .A (nx8894)) ;
    latchr i7_r8_lat_q_3__u1 (.QB (nx8897), .D (nx9318), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_3__u2 (.Y (DecompressedData1[163]), .A (nx8897)) ;
    buf02 i7_r8_lat_q_3__u3 (.Y (nx6607), .A (nx8897)) ;
    latchr i8_r11_lat_q_3__u1 (.QB (nx8900), .D (nx6108), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_3__u2 (.Y (DecompressedData2[163]), .A (nx8900)) ;
    buf02 i8_r11_lat_q_3__u3 (.Y (nx6609), .A (nx8900)) ;
    latchr i7_r8_lat_q_4__u1 (.QB (nx8903), .D (nx9328), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_4__u2 (.Y (DecompressedData1[164]), .A (nx8903)) ;
    buf02 i7_r8_lat_q_4__u3 (.Y (nx6612), .A (nx8903)) ;
    latchr i8_r11_lat_q_4__u1 (.QB (nx8906), .D (nx6132), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_4__u2 (.Y (DecompressedData2[164]), .A (nx8906)) ;
    buf02 i8_r11_lat_q_4__u3 (.Y (nx6615), .A (nx8906)) ;
    latchr i7_r8_lat_q_5__u1 (.QB (nx8909), .D (nx9334), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_5__u2 (.Y (DecompressedData1[165]), .A (nx8909)) ;
    buf02 i7_r8_lat_q_5__u3 (.Y (nx6619), .A (nx8909)) ;
    latchr i8_r11_lat_q_5__u1 (.QB (nx8912), .D (nx6156), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_5__u2 (.Y (DecompressedData2[165]), .A (nx8912)) ;
    buf02 i8_r11_lat_q_5__u3 (.Y (nx6621), .A (nx8912)) ;
    latchr i7_r8_lat_q_6__u1 (.QB (nx8915), .D (nx9338), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_6__u2 (.Y (DecompressedData1[166]), .A (nx8915)) ;
    buf02 i7_r8_lat_q_6__u3 (.Y (nx6624), .A (nx8915)) ;
    latchr i8_r11_lat_q_6__u1 (.QB (nx8918), .D (nx6180), .CLK (nx9380), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_6__u2 (.Y (DecompressedData2[166]), .A (nx8918)) ;
    buf02 i8_r11_lat_q_6__u3 (.Y (nx6627), .A (nx8918)) ;
    latchr i7_r8_lat_q_7__u1 (.QB (nx8921), .D (nx9342), .CLK (nx6010), .R (
           DecompressedData1[255])) ;
    inv01 i7_r8_lat_q_7__u2 (.Y (DecompressedData1[167]), .A (nx8921)) ;
    buf02 i7_r8_lat_q_7__u3 (.Y (nx6631), .A (nx8921)) ;
    latchr i8_r11_lat_q_7__u1 (.QB (nx8924), .D (nx6204), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_7__u2 (.Y (DecompressedData2[167]), .A (nx8924)) ;
    buf02 i8_r11_lat_q_7__u3 (.Y (nx6633), .A (nx8924)) ;
    latchr i7_r7_lat_q_0__u1 (.QB (nx8927), .D (nx9286), .CLK (nx6220), .R (
           DecompressedData1[255])) ;
    inv01 i7_r7_lat_q_0__u2 (.Y (DecompressedData1[168]), .A (nx8927)) ;
    buf02 i7_r7_lat_q_0__u3 (.Y (nx6636), .A (nx8927)) ;
    latchr i8_r11_lat_q_8__u1 (.QB (nx8930), .D (nx6234), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_8__u2 (.Y (DecompressedData2[168]), .A (nx8930)) ;
    buf02 i8_r11_lat_q_8__u3 (.Y (nx6639), .A (nx8930)) ;
    latchr i7_r7_lat_q_1__u1 (.QB (nx8933), .D (nx9300), .CLK (nx6220), .R (
           DecompressedData1[255])) ;
    inv01 i7_r7_lat_q_1__u2 (.Y (DecompressedData1[169]), .A (nx8933)) ;
    buf02 i7_r7_lat_q_1__u3 (.Y (nx6643), .A (nx8933)) ;
    latchr i8_r11_lat_q_9__u1 (.QB (nx8936), .D (nx6258), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_9__u2 (.Y (DecompressedData2[169]), .A (nx8936)) ;
    buf02 i8_r11_lat_q_9__u3 (.Y (nx6645), .A (nx8936)) ;
    latchr i7_r7_lat_q_2__u1 (.QB (nx8939), .D (nx9310), .CLK (nx6220), .R (
           DecompressedData1[255])) ;
    inv01 i7_r7_lat_q_2__u2 (.Y (DecompressedData1[170]), .A (nx8939)) ;
    buf02 i7_r7_lat_q_2__u3 (.Y (nx6648), .A (nx8939)) ;
    latchr i8_r11_lat_q_10__u1 (.QB (nx8942), .D (nx6282), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_10__u2 (.Y (DecompressedData2[170]), .A (nx8942)) ;
    buf02 i8_r11_lat_q_10__u3 (.Y (nx6651), .A (nx8942)) ;
    latchr i7_r7_lat_q_3__u1 (.QB (nx8945), .D (nx9320), .CLK (nx6220), .R (
           DecompressedData1[255])) ;
    inv01 i7_r7_lat_q_3__u2 (.Y (DecompressedData1[171]), .A (nx8945)) ;
    buf02 i7_r7_lat_q_3__u3 (.Y (nx6655), .A (nx8945)) ;
    latchr i8_r11_lat_q_11__u1 (.QB (nx8948), .D (nx6306), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_11__u2 (.Y (DecompressedData2[171]), .A (nx8948)) ;
    buf02 i8_r11_lat_q_11__u3 (.Y (nx6657), .A (nx8948)) ;
    latchr i7_r7_lat_q_4__u1 (.QB (nx8951), .D (nx9330), .CLK (nx6220), .R (
           DecompressedData1[255])) ;
    inv01 i7_r7_lat_q_4__u2 (.Y (DecompressedData1[172]), .A (nx8951)) ;
    buf02 i7_r7_lat_q_4__u3 (.Y (nx6660), .A (nx8951)) ;
    latchr i8_r11_lat_q_12__u1 (.QB (nx8954), .D (nx6330), .CLK (nx9382), .R (
           DecompressedData1[255])) ;
    inv01 i8_r11_lat_q_12__u2 (.Y (DecompressedData2[172]), .A (nx8954)) ;
    buf02 i8_r11_lat_q_12__u3 (.Y (nx6663), .A (nx8954)) ;
    latchr i7_r6_lat_q_0__u1 (.QB (nx8957), .D (nx9286), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_0__u2 (.Y (DecompressedData1[176]), .A (nx8957)) ;
    buf02 i7_r6_lat_q_0__u3 (.Y (nx6679), .A (nx8957)) ;
    latchr i8_r12_lat_q_0__u1 (.QB (nx8960), .D (nx6420), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_0__u2 (.Y (DecompressedData2[176]), .A (nx8960)) ;
    buf02 i8_r12_lat_q_0__u3 (.Y (nx6681), .A (nx8960)) ;
    latchr i7_r6_lat_q_1__u1 (.QB (nx8963), .D (nx9300), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_1__u2 (.Y (DecompressedData1[177]), .A (nx8963)) ;
    buf02 i7_r6_lat_q_1__u3 (.Y (nx6684), .A (nx8963)) ;
    latchr i8_r12_lat_q_1__u1 (.QB (nx8966), .D (nx6444), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_1__u2 (.Y (DecompressedData2[177]), .A (nx8966)) ;
    buf02 i8_r12_lat_q_1__u3 (.Y (nx6687), .A (nx8966)) ;
    latchr i7_r6_lat_q_2__u1 (.QB (nx8969), .D (nx9310), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_2__u2 (.Y (DecompressedData1[178]), .A (nx8969)) ;
    buf02 i7_r6_lat_q_2__u3 (.Y (nx6691), .A (nx8969)) ;
    latchr i8_r12_lat_q_2__u1 (.QB (nx8972), .D (nx6468), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_2__u2 (.Y (DecompressedData2[178]), .A (nx8972)) ;
    buf02 i8_r12_lat_q_2__u3 (.Y (nx6693), .A (nx8972)) ;
    latchr i7_r6_lat_q_3__u1 (.QB (nx8975), .D (nx9320), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_3__u2 (.Y (DecompressedData1[179]), .A (nx8975)) ;
    buf02 i7_r6_lat_q_3__u3 (.Y (nx6696), .A (nx8975)) ;
    latchr i8_r12_lat_q_3__u1 (.QB (nx8978), .D (nx6492), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_3__u2 (.Y (DecompressedData2[179]), .A (nx8978)) ;
    buf02 i8_r12_lat_q_3__u3 (.Y (nx6699), .A (nx8978)) ;
    latchr i7_r6_lat_q_4__u1 (.QB (nx8981), .D (nx9330), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_4__u2 (.Y (DecompressedData1[180]), .A (nx8981)) ;
    buf02 i7_r6_lat_q_4__u3 (.Y (nx6703), .A (nx8981)) ;
    latchr i8_r12_lat_q_4__u1 (.QB (nx8984), .D (nx6516), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_4__u2 (.Y (DecompressedData2[180]), .A (nx8984)) ;
    buf02 i8_r12_lat_q_4__u3 (.Y (nx6705), .A (nx8984)) ;
    latchr i7_r6_lat_q_5__u1 (.QB (nx8987), .D (nx9334), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_5__u2 (.Y (DecompressedData1[181]), .A (nx8987)) ;
    buf02 i7_r6_lat_q_5__u3 (.Y (nx6708), .A (nx8987)) ;
    latchr i8_r12_lat_q_5__u1 (.QB (nx8990), .D (nx6540), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_5__u2 (.Y (DecompressedData2[181]), .A (nx8990)) ;
    buf02 i8_r12_lat_q_5__u3 (.Y (nx6711), .A (nx8990)) ;
    latchr i7_r6_lat_q_6__u1 (.QB (nx8993), .D (nx9338), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_6__u2 (.Y (DecompressedData1[182]), .A (nx8993)) ;
    buf02 i7_r6_lat_q_6__u3 (.Y (nx6715), .A (nx8993)) ;
    latchr i8_r12_lat_q_6__u1 (.QB (nx8996), .D (nx6564), .CLK (nx9384), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_6__u2 (.Y (DecompressedData2[182]), .A (nx8996)) ;
    buf02 i8_r12_lat_q_6__u3 (.Y (nx6717), .A (nx8996)) ;
    latchr i7_r6_lat_q_7__u1 (.QB (nx8999), .D (nx9342), .CLK (nx6394), .R (
           DecompressedData1[255])) ;
    inv01 i7_r6_lat_q_7__u2 (.Y (DecompressedData1[183]), .A (nx8999)) ;
    buf02 i7_r6_lat_q_7__u3 (.Y (nx6720), .A (nx8999)) ;
    latchr i8_r12_lat_q_7__u1 (.QB (nx9002), .D (nx6588), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_7__u2 (.Y (DecompressedData2[183]), .A (nx9002)) ;
    buf02 i8_r12_lat_q_7__u3 (.Y (nx6723), .A (nx9002)) ;
    latchr i7_r5_lat_q_0__u1 (.QB (nx9005), .D (nx9286), .CLK (nx6604), .R (
           DecompressedData1[255])) ;
    inv01 i7_r5_lat_q_0__u2 (.Y (DecompressedData1[184]), .A (nx9005)) ;
    buf02 i7_r5_lat_q_0__u3 (.Y (nx6727), .A (nx9005)) ;
    latchr i8_r12_lat_q_8__u1 (.QB (nx9008), .D (nx6618), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_8__u2 (.Y (DecompressedData2[184]), .A (nx9008)) ;
    buf02 i8_r12_lat_q_8__u3 (.Y (nx6729), .A (nx9008)) ;
    latchr i7_r5_lat_q_1__u1 (.QB (nx9011), .D (nx9300), .CLK (nx6604), .R (
           DecompressedData1[255])) ;
    inv01 i7_r5_lat_q_1__u2 (.Y (DecompressedData1[185]), .A (nx9011)) ;
    buf02 i7_r5_lat_q_1__u3 (.Y (nx6732), .A (nx9011)) ;
    latchr i8_r12_lat_q_9__u1 (.QB (nx9014), .D (nx6642), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_9__u2 (.Y (DecompressedData2[185]), .A (nx9014)) ;
    buf02 i8_r12_lat_q_9__u3 (.Y (nx6734), .A (nx9014)) ;
    latchr i7_r5_lat_q_2__u1 (.QB (nx9017), .D (nx9310), .CLK (nx6604), .R (
           DecompressedData1[255])) ;
    inv01 i7_r5_lat_q_2__u2 (.Y (DecompressedData1[186]), .A (nx9017)) ;
    buf02 i7_r5_lat_q_2__u3 (.Y (nx6737), .A (nx9017)) ;
    latchr i8_r12_lat_q_10__u1 (.QB (nx9020), .D (nx6666), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_10__u2 (.Y (DecompressedData2[186]), .A (nx9020)) ;
    buf02 i8_r12_lat_q_10__u3 (.Y (nx6739), .A (nx9020)) ;
    latchr i7_r5_lat_q_3__u1 (.QB (nx9023), .D (nx9320), .CLK (nx6604), .R (
           DecompressedData1[255])) ;
    inv01 i7_r5_lat_q_3__u2 (.Y (DecompressedData1[187]), .A (nx9023)) ;
    buf02 i7_r5_lat_q_3__u3 (.Y (nx6742), .A (nx9023)) ;
    latchr i8_r12_lat_q_11__u1 (.QB (nx9026), .D (nx6690), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_11__u2 (.Y (DecompressedData2[187]), .A (nx9026)) ;
    buf02 i8_r12_lat_q_11__u3 (.Y (nx6744), .A (nx9026)) ;
    latchr i7_r5_lat_q_4__u1 (.QB (nx9029), .D (nx9330), .CLK (nx6604), .R (
           DecompressedData1[255])) ;
    inv01 i7_r5_lat_q_4__u2 (.Y (DecompressedData1[188]), .A (nx9029)) ;
    buf02 i7_r5_lat_q_4__u3 (.Y (nx6747), .A (nx9029)) ;
    latchr i8_r12_lat_q_12__u1 (.QB (nx9032), .D (nx6714), .CLK (nx9386), .R (
           DecompressedData1[255])) ;
    inv01 i8_r12_lat_q_12__u2 (.Y (DecompressedData2[188]), .A (nx9032)) ;
    buf02 i8_r12_lat_q_12__u3 (.Y (nx6749), .A (nx9032)) ;
    latchr i7_r4_lat_q_0__u1 (.QB (nx9035), .D (nx9286), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_0__u2 (.Y (DecompressedData1[192]), .A (nx9035)) ;
    buf02 i7_r4_lat_q_0__u3 (.Y (nx6764), .A (nx9035)) ;
    latchr i8_r13_lat_q_0__u1 (.QB (nx9038), .D (nx6812), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_0__u2 (.Y (DecompressedData2[192]), .A (nx9038)) ;
    buf02 i8_r13_lat_q_0__u3 (.Y (nx6766), .A (nx9038)) ;
    latchr i7_r4_lat_q_1__u1 (.QB (nx9041), .D (nx9300), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_1__u2 (.Y (DecompressedData1[193]), .A (nx9041)) ;
    buf02 i7_r4_lat_q_1__u3 (.Y (nx6769), .A (nx9041)) ;
    latchr i8_r13_lat_q_1__u1 (.QB (nx9044), .D (nx6836), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_1__u2 (.Y (DecompressedData2[193]), .A (nx9044)) ;
    buf02 i8_r13_lat_q_1__u3 (.Y (nx6771), .A (nx9044)) ;
    latchr i7_r4_lat_q_2__u1 (.QB (nx9047), .D (nx9310), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_2__u2 (.Y (DecompressedData1[194]), .A (nx9047)) ;
    buf02 i7_r4_lat_q_2__u3 (.Y (nx6775), .A (nx9047)) ;
    latchr i8_r13_lat_q_2__u1 (.QB (nx9050), .D (nx6860), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_2__u2 (.Y (DecompressedData2[194]), .A (nx9050)) ;
    buf02 i8_r13_lat_q_2__u3 (.Y (nx6777), .A (nx9050)) ;
    latchr i7_r4_lat_q_3__u1 (.QB (nx9053), .D (nx9320), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_3__u2 (.Y (DecompressedData1[195]), .A (nx9053)) ;
    buf02 i7_r4_lat_q_3__u3 (.Y (nx6781), .A (nx9053)) ;
    latchr i8_r13_lat_q_3__u1 (.QB (nx9056), .D (nx6884), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_3__u2 (.Y (DecompressedData2[195]), .A (nx9056)) ;
    buf02 i8_r13_lat_q_3__u3 (.Y (nx6783), .A (nx9056)) ;
    latchr i7_r4_lat_q_4__u1 (.QB (nx9059), .D (nx9330), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_4__u2 (.Y (DecompressedData1[196]), .A (nx9059)) ;
    buf02 i7_r4_lat_q_4__u3 (.Y (nx6787), .A (nx9059)) ;
    latchr i8_r13_lat_q_4__u1 (.QB (nx9062), .D (nx6908), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_4__u2 (.Y (DecompressedData2[196]), .A (nx9062)) ;
    buf02 i8_r13_lat_q_4__u3 (.Y (nx6789), .A (nx9062)) ;
    latchr i7_r4_lat_q_5__u1 (.QB (nx9065), .D (nx9334), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_5__u2 (.Y (DecompressedData1[197]), .A (nx9065)) ;
    buf02 i7_r4_lat_q_5__u3 (.Y (nx6792), .A (nx9065)) ;
    latchr i8_r13_lat_q_5__u1 (.QB (nx9068), .D (nx6932), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_5__u2 (.Y (DecompressedData2[197]), .A (nx9068)) ;
    buf02 i8_r13_lat_q_5__u3 (.Y (nx6794), .A (nx9068)) ;
    latchr i7_r4_lat_q_6__u1 (.QB (nx9071), .D (nx9338), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_6__u2 (.Y (DecompressedData1[198]), .A (nx9071)) ;
    buf02 i7_r4_lat_q_6__u3 (.Y (nx6797), .A (nx9071)) ;
    latchr i8_r13_lat_q_6__u1 (.QB (nx9074), .D (nx6956), .CLK (nx9388), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_6__u2 (.Y (DecompressedData2[198]), .A (nx9074)) ;
    buf02 i8_r13_lat_q_6__u3 (.Y (nx6799), .A (nx9074)) ;
    latchr i7_r4_lat_q_7__u1 (.QB (nx9077), .D (nx9342), .CLK (nx6786), .R (
           DecompressedData1[255])) ;
    inv01 i7_r4_lat_q_7__u2 (.Y (DecompressedData1[199]), .A (nx9077)) ;
    buf02 i7_r4_lat_q_7__u3 (.Y (nx6803), .A (nx9077)) ;
    latchr i8_r13_lat_q_7__u1 (.QB (nx9080), .D (nx6980), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_7__u2 (.Y (DecompressedData2[199]), .A (nx9080)) ;
    buf02 i8_r13_lat_q_7__u3 (.Y (nx6805), .A (nx9080)) ;
    latchr i7_r3_lat_q_0__u1 (.QB (nx9083), .D (nx9286), .CLK (nx6996), .R (
           DecompressedData1[255])) ;
    inv01 i7_r3_lat_q_0__u2 (.Y (DecompressedData1[200]), .A (nx9083)) ;
    buf02 i7_r3_lat_q_0__u3 (.Y (nx6809), .A (nx9083)) ;
    latchr i8_r13_lat_q_8__u1 (.QB (nx9086), .D (nx7010), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_8__u2 (.Y (DecompressedData2[200]), .A (nx9086)) ;
    buf02 i8_r13_lat_q_8__u3 (.Y (nx6811), .A (nx9086)) ;
    latchr i7_r3_lat_q_1__u1 (.QB (nx9089), .D (nx9300), .CLK (nx6996), .R (
           DecompressedData1[255])) ;
    inv01 i7_r3_lat_q_1__u2 (.Y (DecompressedData1[201]), .A (nx9089)) ;
    buf02 i7_r3_lat_q_1__u3 (.Y (nx6815), .A (nx9089)) ;
    latchr i8_r13_lat_q_9__u1 (.QB (nx9092), .D (nx7034), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_9__u2 (.Y (DecompressedData2[201]), .A (nx9092)) ;
    buf02 i8_r13_lat_q_9__u3 (.Y (nx6817), .A (nx9092)) ;
    latchr i7_r3_lat_q_2__u1 (.QB (nx9095), .D (nx9310), .CLK (nx6996), .R (
           DecompressedData1[255])) ;
    inv01 i7_r3_lat_q_2__u2 (.Y (DecompressedData1[202]), .A (nx9095)) ;
    buf02 i7_r3_lat_q_2__u3 (.Y (nx6821), .A (nx9095)) ;
    latchr i8_r13_lat_q_10__u1 (.QB (nx9098), .D (nx7058), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_10__u2 (.Y (DecompressedData2[202]), .A (nx9098)) ;
    buf02 i8_r13_lat_q_10__u3 (.Y (nx6823), .A (nx9098)) ;
    latchr i7_r3_lat_q_3__u1 (.QB (nx9101), .D (nx9320), .CLK (nx6996), .R (
           DecompressedData1[255])) ;
    inv01 i7_r3_lat_q_3__u2 (.Y (DecompressedData1[203]), .A (nx9101)) ;
    buf02 i7_r3_lat_q_3__u3 (.Y (nx6826), .A (nx9101)) ;
    latchr i8_r13_lat_q_11__u1 (.QB (nx9104), .D (nx7082), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_11__u2 (.Y (DecompressedData2[203]), .A (nx9104)) ;
    buf02 i8_r13_lat_q_11__u3 (.Y (nx6828), .A (nx9104)) ;
    latchr i7_r3_lat_q_4__u1 (.QB (nx9107), .D (nx9330), .CLK (nx6996), .R (
           DecompressedData1[255])) ;
    inv01 i7_r3_lat_q_4__u2 (.Y (DecompressedData1[204]), .A (nx9107)) ;
    buf02 i7_r3_lat_q_4__u3 (.Y (nx6831), .A (nx9107)) ;
    latchr i8_r13_lat_q_12__u1 (.QB (nx9110), .D (nx7106), .CLK (nx9390), .R (
           DecompressedData1[255])) ;
    inv01 i8_r13_lat_q_12__u2 (.Y (DecompressedData2[204]), .A (nx9110)) ;
    buf02 i8_r13_lat_q_12__u3 (.Y (nx6833), .A (nx9110)) ;
    latchr i7_r2_lat_q_0__u1 (.QB (nx9113), .D (nx9286), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_0__u2 (.Y (DecompressedData1[208]), .A (nx9113)) ;
    buf02 i7_r2_lat_q_0__u3 (.Y (nx6849), .A (nx9113)) ;
    latchr i8_r14_lat_q_0__u1 (.QB (nx9116), .D (nx7196), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_0__u2 (.Y (DecompressedData2[208]), .A (nx9116)) ;
    buf02 i8_r14_lat_q_0__u3 (.Y (nx6851), .A (nx9116)) ;
    latchr i7_r2_lat_q_1__u1 (.QB (nx9119), .D (nx9300), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_1__u2 (.Y (DecompressedData1[209]), .A (nx9119)) ;
    buf02 i7_r2_lat_q_1__u3 (.Y (nx6854), .A (nx9119)) ;
    latchr i8_r14_lat_q_1__u1 (.QB (nx9122), .D (nx7220), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_1__u2 (.Y (DecompressedData2[209]), .A (nx9122)) ;
    buf02 i8_r14_lat_q_1__u3 (.Y (nx6857), .A (nx9122)) ;
    latchr i7_r2_lat_q_2__u1 (.QB (nx9125), .D (nx9310), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_2__u2 (.Y (DecompressedData1[210]), .A (nx9125)) ;
    buf02 i7_r2_lat_q_2__u3 (.Y (nx6861), .A (nx9125)) ;
    latchr i8_r14_lat_q_2__u1 (.QB (nx9128), .D (nx7244), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_2__u2 (.Y (DecompressedData2[210]), .A (nx9128)) ;
    buf02 i8_r14_lat_q_2__u3 (.Y (nx6863), .A (nx9128)) ;
    latchr i7_r2_lat_q_3__u1 (.QB (nx9131), .D (nx9320), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_3__u2 (.Y (DecompressedData1[211]), .A (nx9131)) ;
    buf02 i7_r2_lat_q_3__u3 (.Y (nx6866), .A (nx9131)) ;
    latchr i8_r14_lat_q_3__u1 (.QB (nx9134), .D (nx7268), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_3__u2 (.Y (DecompressedData2[211]), .A (nx9134)) ;
    buf02 i8_r14_lat_q_3__u3 (.Y (nx6869), .A (nx9134)) ;
    latchr i7_r2_lat_q_4__u1 (.QB (nx9137), .D (nx9330), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_4__u2 (.Y (DecompressedData1[212]), .A (nx9137)) ;
    buf02 i7_r2_lat_q_4__u3 (.Y (nx6873), .A (nx9137)) ;
    latchr i8_r14_lat_q_4__u1 (.QB (nx9140), .D (nx7292), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_4__u2 (.Y (DecompressedData2[212]), .A (nx9140)) ;
    buf02 i8_r14_lat_q_4__u3 (.Y (nx6875), .A (nx9140)) ;
    latchr i7_r2_lat_q_5__u1 (.QB (nx9143), .D (nx9334), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_5__u2 (.Y (DecompressedData1[213]), .A (nx9143)) ;
    buf02 i7_r2_lat_q_5__u3 (.Y (nx6878), .A (nx9143)) ;
    latchr i8_r14_lat_q_5__u1 (.QB (nx9146), .D (nx7316), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_5__u2 (.Y (DecompressedData2[213]), .A (nx9146)) ;
    buf02 i8_r14_lat_q_5__u3 (.Y (nx6881), .A (nx9146)) ;
    latchr i7_r2_lat_q_6__u1 (.QB (nx9149), .D (nx9338), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_6__u2 (.Y (DecompressedData1[214]), .A (nx9149)) ;
    buf02 i7_r2_lat_q_6__u3 (.Y (nx6885), .A (nx9149)) ;
    latchr i8_r14_lat_q_6__u1 (.QB (nx9152), .D (nx7340), .CLK (nx9392), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_6__u2 (.Y (DecompressedData2[214]), .A (nx9152)) ;
    buf02 i8_r14_lat_q_6__u3 (.Y (nx6887), .A (nx9152)) ;
    latchr i7_r2_lat_q_7__u1 (.QB (nx9155), .D (nx9342), .CLK (nx7170), .R (
           DecompressedData1[255])) ;
    inv01 i7_r2_lat_q_7__u2 (.Y (DecompressedData1[215]), .A (nx9155)) ;
    buf02 i7_r2_lat_q_7__u3 (.Y (nx6890), .A (nx9155)) ;
    latchr i8_r14_lat_q_7__u1 (.QB (nx9158), .D (nx7364), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_7__u2 (.Y (DecompressedData2[215]), .A (nx9158)) ;
    buf02 i8_r14_lat_q_7__u3 (.Y (nx6893), .A (nx9158)) ;
    latchr i7_r1_lat_q_0__u1 (.QB (nx9161), .D (nx9286), .CLK (nx7380), .R (
           DecompressedData1[255])) ;
    inv01 i7_r1_lat_q_0__u2 (.Y (DecompressedData1[216]), .A (nx9161)) ;
    buf02 i7_r1_lat_q_0__u3 (.Y (nx6897), .A (nx9161)) ;
    latchr i8_r14_lat_q_8__u1 (.QB (nx9164), .D (nx7394), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_8__u2 (.Y (DecompressedData2[216]), .A (nx9164)) ;
    buf02 i8_r14_lat_q_8__u3 (.Y (nx6899), .A (nx9164)) ;
    latchr i7_r1_lat_q_1__u1 (.QB (nx9167), .D (nx9300), .CLK (nx7380), .R (
           DecompressedData1[255])) ;
    inv01 i7_r1_lat_q_1__u2 (.Y (DecompressedData1[217]), .A (nx9167)) ;
    buf02 i7_r1_lat_q_1__u3 (.Y (nx6902), .A (nx9167)) ;
    latchr i8_r14_lat_q_9__u1 (.QB (nx9170), .D (nx7418), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_9__u2 (.Y (DecompressedData2[217]), .A (nx9170)) ;
    buf02 i8_r14_lat_q_9__u3 (.Y (nx6905), .A (nx9170)) ;
    latchr i7_r1_lat_q_2__u1 (.QB (nx9173), .D (nx9310), .CLK (nx7380), .R (
           DecompressedData1[255])) ;
    inv01 i7_r1_lat_q_2__u2 (.Y (DecompressedData1[218]), .A (nx9173)) ;
    buf02 i7_r1_lat_q_2__u3 (.Y (nx6909), .A (nx9173)) ;
    latchr i8_r14_lat_q_10__u1 (.QB (nx9176), .D (nx7442), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_10__u2 (.Y (DecompressedData2[218]), .A (nx9176)) ;
    buf02 i8_r14_lat_q_10__u3 (.Y (nx6911), .A (nx9176)) ;
    latchr i7_r1_lat_q_3__u1 (.QB (nx9179), .D (nx9320), .CLK (nx7380), .R (
           DecompressedData1[255])) ;
    inv01 i7_r1_lat_q_3__u2 (.Y (DecompressedData1[219]), .A (nx9179)) ;
    buf02 i7_r1_lat_q_3__u3 (.Y (nx6914), .A (nx9179)) ;
    latchr i8_r14_lat_q_11__u1 (.QB (nx9182), .D (nx7466), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_11__u2 (.Y (DecompressedData2[219]), .A (nx9182)) ;
    buf02 i8_r14_lat_q_11__u3 (.Y (nx6917), .A (nx9182)) ;
    latchr i7_r1_lat_q_4__u1 (.QB (nx9185), .D (nx9330), .CLK (nx7380), .R (
           DecompressedData1[255])) ;
    inv01 i7_r1_lat_q_4__u2 (.Y (DecompressedData1[220]), .A (nx9185)) ;
    buf02 i7_r1_lat_q_4__u3 (.Y (nx6921), .A (nx9185)) ;
    latchr i8_r14_lat_q_12__u1 (.QB (nx9188), .D (nx7490), .CLK (nx9394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r14_lat_q_12__u2 (.Y (DecompressedData2[220]), .A (nx9188)) ;
    buf02 i8_r14_lat_q_12__u3 (.Y (nx6923), .A (nx9188)) ;
    latchr i8_r15_lat_q_0__u1 (.QB (nx9191), .D (nx1192), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_0__u2 (.Y (DecompressedData2[224]), .A (nx9191)) ;
    buf02 i8_r15_lat_q_0__u3 (.Y (nx6939), .A (nx9191)) ;
    latchr i8_r15_lat_q_1__u1 (.QB (nx9194), .D (nx1206), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_1__u2 (.Y (DecompressedData2[225]), .A (nx9194)) ;
    buf02 i8_r15_lat_q_1__u3 (.Y (nx6943), .A (nx9194)) ;
    latchr i8_r15_lat_q_2__u1 (.QB (nx9197), .D (nx1220), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_2__u2 (.Y (DecompressedData2[226]), .A (nx9197)) ;
    buf02 i8_r15_lat_q_2__u3 (.Y (nx6946), .A (nx9197)) ;
    latchr i8_r15_lat_q_3__u1 (.QB (nx9200), .D (nx1234), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_3__u2 (.Y (DecompressedData2[227]), .A (nx9200)) ;
    buf02 i8_r15_lat_q_3__u3 (.Y (nx6949), .A (nx9200)) ;
    latchr i8_r15_lat_q_4__u1 (.QB (nx9203), .D (nx1248), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_4__u2 (.Y (DecompressedData2[228]), .A (nx9203)) ;
    buf02 i8_r15_lat_q_4__u3 (.Y (nx6953), .A (nx9203)) ;
    latchr i8_r15_lat_q_5__u1 (.QB (nx9206), .D (nx1262), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_5__u2 (.Y (DecompressedData2[229]), .A (nx9206)) ;
    buf02 i8_r15_lat_q_5__u3 (.Y (nx6957), .A (nx9206)) ;
    latchr i8_r15_lat_q_6__u1 (.QB (nx9209), .D (nx1276), .CLK (nx9274), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_6__u2 (.Y (DecompressedData2[230]), .A (nx9209)) ;
    buf02 i8_r15_lat_q_6__u3 (.Y (nx6960), .A (nx9209)) ;
    latchr i8_r15_lat_q_7__u1 (.QB (nx9212), .D (nx1290), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_7__u2 (.Y (DecompressedData2[231]), .A (nx9212)) ;
    buf02 i8_r15_lat_q_7__u3 (.Y (nx6963), .A (nx9212)) ;
    latchr i8_r15_lat_q_8__u1 (.QB (nx9215), .D (nx1304), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_8__u2 (.Y (DecompressedData2[232]), .A (nx9215)) ;
    buf02 i8_r15_lat_q_8__u3 (.Y (nx6967), .A (nx9215)) ;
    latchr i8_r15_lat_q_9__u1 (.QB (nx9218), .D (nx1318), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_9__u2 (.Y (DecompressedData2[233]), .A (nx9218)) ;
    buf02 i8_r15_lat_q_9__u3 (.Y (nx6970), .A (nx9218)) ;
    latchr i8_r15_lat_q_10__u1 (.QB (nx9221), .D (nx1332), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_10__u2 (.Y (DecompressedData2[234]), .A (nx9221)) ;
    buf02 i8_r15_lat_q_10__u3 (.Y (nx6973), .A (nx9221)) ;
    latchr i8_r15_lat_q_11__u1 (.QB (nx9224), .D (nx1346), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_11__u2 (.Y (DecompressedData2[235]), .A (nx9224)) ;
    buf02 i8_r15_lat_q_11__u3 (.Y (nx6977), .A (nx9224)) ;
    latchr i8_r15_lat_q_12__u1 (.QB (nx9227), .D (nx1360), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_12__u2 (.Y (DecompressedData2[236]), .A (nx9227)) ;
    buf02 i8_r15_lat_q_12__u3 (.Y (nx6981), .A (nx9227)) ;
    latchr i8_r15_lat_q_13__u1 (.QB (nx9230), .D (nx1374), .CLK (nx1186), .R (
           DecompressedData1[255])) ;
    inv01 i8_r15_lat_q_13__u2 (.Y (DecompressedData2[239]), .A (nx9230)) ;
    buf02 i8_r15_lat_q_13__u3 (.Y (nx6984), .A (nx9230)) ;
    latchr i8_r16_lat_q_0__u1 (.QB (nx9233), .D (nx1398), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_0__u2 (.Y (DecompressedData2[240]), .A (nx9233)) ;
    buf02 i8_r16_lat_q_0__u3 (.Y (nx6987), .A (nx9233)) ;
    latchr i8_r16_lat_q_1__u1 (.QB (nx9236), .D (nx1410), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_1__u2 (.Y (DecompressedData2[241]), .A (nx9236)) ;
    buf02 i8_r16_lat_q_1__u3 (.Y (nx6991), .A (nx9236)) ;
    latchr i8_r16_lat_q_2__u1 (.QB (nx9239), .D (nx1422), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_2__u2 (.Y (DecompressedData2[242]), .A (nx9239)) ;
    buf02 i8_r16_lat_q_2__u3 (.Y (nx6995), .A (nx9239)) ;
    latchr i8_r16_lat_q_3__u1 (.QB (nx9242), .D (nx1434), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_3__u2 (.Y (DecompressedData2[243]), .A (nx9242)) ;
    buf02 i8_r16_lat_q_3__u3 (.Y (nx6999), .A (nx9242)) ;
    latchr i8_r16_lat_q_4__u1 (.QB (nx9245), .D (nx1446), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_4__u2 (.Y (DecompressedData2[244]), .A (nx9245)) ;
    buf02 i8_r16_lat_q_4__u3 (.Y (nx7002), .A (nx9245)) ;
    latchr i8_r16_lat_q_5__u1 (.QB (nx9248), .D (nx1458), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_5__u2 (.Y (DecompressedData2[245]), .A (nx9248)) ;
    buf02 i8_r16_lat_q_5__u3 (.Y (nx7005), .A (nx9248)) ;
    latchr i8_r16_lat_q_6__u1 (.QB (nx9251), .D (nx1470), .CLK (nx9276), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_6__u2 (.Y (DecompressedData2[246]), .A (nx9251)) ;
    buf02 i8_r16_lat_q_6__u3 (.Y (nx7009), .A (nx9251)) ;
    latchr i8_r16_lat_q_7__u1 (.QB (nx9254), .D (nx1482), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_7__u2 (.Y (DecompressedData2[247]), .A (nx9254)) ;
    buf02 i8_r16_lat_q_7__u3 (.Y (nx7013), .A (nx9254)) ;
    latchr i8_r16_lat_q_8__u1 (.QB (nx9257), .D (nx1494), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_8__u2 (.Y (DecompressedData2[248]), .A (nx9257)) ;
    buf02 i8_r16_lat_q_8__u3 (.Y (nx7016), .A (nx9257)) ;
    latchr i8_r16_lat_q_9__u1 (.QB (nx9260), .D (nx1506), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_9__u2 (.Y (DecompressedData2[249]), .A (nx9260)) ;
    buf02 i8_r16_lat_q_9__u3 (.Y (nx7019), .A (nx9260)) ;
    latchr i8_r16_lat_q_10__u1 (.QB (nx9263), .D (nx1518), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_10__u2 (.Y (DecompressedData2[250]), .A (nx9263)) ;
    buf02 i8_r16_lat_q_10__u3 (.Y (nx7023), .A (nx9263)) ;
    latchr i8_r16_lat_q_11__u1 (.QB (nx9266), .D (nx1530), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_11__u2 (.Y (DecompressedData2[251]), .A (nx9266)) ;
    buf02 i8_r16_lat_q_11__u3 (.Y (nx7026), .A (nx9266)) ;
    latchr i8_r16_lat_q_12__u1 (.QB (nx9269), .D (nx1542), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_12__u2 (.Y (DecompressedData2[252]), .A (nx9269)) ;
    buf02 i8_r16_lat_q_12__u3 (.Y (nx7029), .A (nx9269)) ;
    latchr i8_r16_lat_q_13__u1 (.QB (nx9272), .D (nx1554), .CLK (nx1394), .R (
           DecompressedData1[255])) ;
    inv01 i8_r16_lat_q_13__u2 (.Y (DecompressedData2[255]), .A (nx9272)) ;
    buf02 i8_r16_lat_q_13__u3 (.Y (nx7033), .A (nx9272)) ;
    nand02 ix9273 (.Y (nx9274), .A0 (nx5212), .A1 (nx5215)) ;
    nand02 ix9275 (.Y (nx9276), .A0 (nx5266), .A1 (nx5259)) ;
    inv01 ix9277 (.Y (nx9278), .A (nx2086)) ;
    inv02 ix9279 (.Y (nx9280), .A (nx9278)) ;
    inv02 ix9281 (.Y (nx9282), .A (nx9278)) ;
    inv02 ix9283 (.Y (nx9284), .A (nx9278)) ;
    inv02 ix9285 (.Y (nx9286), .A (nx9278)) ;
    inv02 ix9287 (.Y (nx9288), .A (nx7539)) ;
    inv02 ix9289 (.Y (nx9290), .A (nx7539)) ;
    inv01 ix9291 (.Y (nx9292), .A (nx2134)) ;
    inv02 ix9293 (.Y (nx9294), .A (nx9292)) ;
    inv02 ix9295 (.Y (nx9296), .A (nx9292)) ;
    inv02 ix9297 (.Y (nx9298), .A (nx9292)) ;
    inv02 ix9299 (.Y (nx9300), .A (nx9292)) ;
    inv01 ix9301 (.Y (nx9302), .A (nx2160)) ;
    inv02 ix9303 (.Y (nx9304), .A (nx9302)) ;
    inv02 ix9305 (.Y (nx9306), .A (nx9302)) ;
    inv02 ix9307 (.Y (nx9308), .A (nx9302)) ;
    inv02 ix9309 (.Y (nx9310), .A (nx9302)) ;
    inv01 ix9311 (.Y (nx9312), .A (nx2186)) ;
    inv02 ix9313 (.Y (nx9314), .A (nx9312)) ;
    inv02 ix9315 (.Y (nx9316), .A (nx9312)) ;
    inv02 ix9317 (.Y (nx9318), .A (nx9312)) ;
    inv02 ix9319 (.Y (nx9320), .A (nx9312)) ;
    inv01 ix9321 (.Y (nx9322), .A (nx2212)) ;
    inv02 ix9323 (.Y (nx9324), .A (nx9322)) ;
    inv02 ix9325 (.Y (nx9326), .A (nx9322)) ;
    inv02 ix9327 (.Y (nx9328), .A (nx9322)) ;
    inv02 ix9329 (.Y (nx9330), .A (nx9322)) ;
    inv02 ix9331 (.Y (nx9332), .A (nx7551)) ;
    inv02 ix9333 (.Y (nx9334), .A (nx7551)) ;
    inv02 ix9335 (.Y (nx9336), .A (nx7557)) ;
    inv02 ix9337 (.Y (nx9338), .A (nx7557)) ;
    inv02 ix9339 (.Y (nx9340), .A (nx7563)) ;
    inv02 ix9341 (.Y (nx9342), .A (nx7563)) ;
    inv02 ix9343 (.Y (nx9344), .A (nx7577)) ;
    inv02 ix9345 (.Y (nx9346), .A (nx7577)) ;
    inv02 ix9347 (.Y (nx9348), .A (nx7589)) ;
    inv02 ix9349 (.Y (nx9350), .A (nx7589)) ;
    inv02 ix9351 (.Y (nx9352), .A (nx7601)) ;
    inv02 ix9353 (.Y (nx9354), .A (nx7601)) ;
    inv02 ix9355 (.Y (nx9356), .A (nx7613)) ;
    inv02 ix9357 (.Y (nx9358), .A (nx7613)) ;
    inv02 ix9359 (.Y (nx9360), .A (nx7625)) ;
    inv02 ix9361 (.Y (nx9362), .A (nx7625)) ;
    inv02 ix9363 (.Y (nx9364), .A (nx7645)) ;
    inv02 ix9365 (.Y (nx9366), .A (nx7645)) ;
    inv02 ix9367 (.Y (nx9368), .A (nx7657)) ;
    inv02 ix9369 (.Y (nx9370), .A (nx7657)) ;
    inv02 ix9371 (.Y (nx9372), .A (nx7669)) ;
    inv02 ix9373 (.Y (nx9374), .A (nx7669)) ;
    inv02 ix9375 (.Y (nx9376), .A (nx7681)) ;
    inv02 ix9377 (.Y (nx9378), .A (nx7681)) ;
    inv02 ix9379 (.Y (nx9380), .A (nx7693)) ;
    inv02 ix9381 (.Y (nx9382), .A (nx7693)) ;
    inv02 ix9383 (.Y (nx9384), .A (nx7705)) ;
    inv02 ix9385 (.Y (nx9386), .A (nx7705)) ;
    inv02 ix9387 (.Y (nx9388), .A (nx7717)) ;
    inv02 ix9389 (.Y (nx9390), .A (nx7717)) ;
    inv02 ix9391 (.Y (nx9392), .A (nx7729)) ;
    inv02 ix9393 (.Y (nx9394), .A (nx7729)) ;
    inv02 ix9395 (.Y (nx9396), .A (nx7401)) ;
    inv02 ix9397 (.Y (nx9398), .A (nx7889)) ;
    inv02 ix9399 (.Y (nx9400), .A (nx7889)) ;
    inv02 ix9401 (.Y (nx9402), .A (nx7889)) ;
    inv02 ix9403 (.Y (nx9404), .A (nx7889)) ;
    inv02 ix9405 (.Y (nx9406), .A (nx7889)) ;
    inv02 ix9407 (.Y (nx9408), .A (nx7889)) ;
endmodule

