
-- 
-- Definition of  IOCHIP
-- 
--      Wed Apr 24 13:15:34 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity IOCHIP is
   port (
      OuterRead : IN std_logic ;
      OuterWrite : IN std_logic ;
      ActivateOuterAddress : IN std_logic ;
      INCEnable : IN std_logic ;
      PDone : IN std_logic ;
      OuterAddress : IN std_logic_vector (15 DOWNTO 0) ;
      ResultIn : IN std_logic_vector (3 DOWNTO 0) ;
      CLK : IN std_logic ;
      LP : IN std_logic ;
      INTR : IN std_logic ;
      CNNIMGLOAD : IN std_logic ;
      Rst : IN std_logic ;
      EnableReadingFromCPU : INOUT std_logic ;
      DecompressionDone : INOUT std_logic ;
      DecompressionDone1 : INOUT std_logic ;
      DecompressionDone2 : INOUT std_logic ;
      readenable : INOUT std_logic ;
      DataBus : IN std_logic_vector (15 DOWNTO 0) ;
      Address : INOUT std_logic_vector (15 DOWNTO 0) ;
      DecompressedData : INOUT std_logic_vector (255 DOWNTO 0) ;
      DecompressedData1 : INOUT std_logic_vector (255 DOWNTO 0) ;
      DecompressedData2 : INOUT std_logic_vector (255 DOWNTO 0) ;
      EnableReadingFromCPU1 : INOUT std_logic ;
      EnableReadingFromCPU2 : INOUT std_logic ;
      loadingimg : INOUT std_logic ;
      loadingCNN : INOUT std_logic ;
      PClk : OUT std_logic ;
      DataFromRam : OUT std_logic_vector (255 DOWNTO 0) ;
      Result : INOUT std_logic_vector (3 DOWNTO 0) ;
      Done : INOUT std_logic ;
      ProcessEnable : OUT std_logic) ;
end IOCHIP ;

architecture arch of IOCHIP is
   signal ProcessEnable_EXMPLR, i8_reset2, nx2, loadenable, nx8, nx14, nx22, 
      nx28, nx32, nx44, nx46, nx52, nx54, nx62, nx66, nx70, nx74, nx82, 
      i8_read2, zed, i8_counterout1_1, i8_reset1, nx98, i8_counterout1_7, 
      nx102, nx104, nx110, i8_counterout1_5, i8_counterout1_4, 
      i8_counterout1_3, i8_counterout1_2, nx3092, i8_counterout1_0, nx128, 
      nx136, nx152, nx3093, nx182, nx3095, nx206, nx3097, nx230, nx3099, 
      nx254, nx268, nx278, nx282, nx298, i8_nx74, nx314, nx316, nx330, nx340, 
      nx356, nx360, nx362, i8_counterout2_5, nx370, nx374, nx376, 
      i8_counterout2_4, nx3100, i8_counterout2_3, nx3101, i8_counterout2_2, 
      nx3102, i8_counterout2_1, i8_counterout2_0, nx396, nx408, nx424, nx444, 
      nx458, nx464, i8_counterout2_7, i8_counterout2_6, nx480, nx494, nx514, 
      nx520, nx528, nx532, nx536, nx3104, nx540, nx546, nx558, nx560, nx572, 
      i8_loadenableD, nx588, nx602, nx610, nx618, nx622, i7_tmp, 
      i7_counterout1_7, i7_start, nx638, i7_reset2, i7_read2, 
      i7_counterout2_7, nx648, nx650, nx654, i7_counterout2_6, 
      i7_counterout2_5, nx3107, i7_counterout2_4, nx3109, i7_counterout2_3, 
      nx3111, i7_counterout2_2, i7_counterout2_1, i7_counterout2_0, nx674, 
      nx690, nx708, nx724, nx740, nx758, nx772, nx796, nx802, nx808, nx812, 
      nx814, NOT_nx814, nx818, nx830, nx836, i7_loadenableD, nx846, nx856, 
      i7_counterout1_6, nx862, nx874, i7_counterout1_5, nx3115, 
      i7_counterout1_4, nx3116, nx894, i7_counterout1_3, nx3117, nx912, 
      i7_counterout1_2, nx3118, nx926, i7_counterout1_1, nx940, 
      i7_counterout1_0, nx952, nx960, nx974, nx994, nx1014, nx1034, nx1054, 
      nx1058, nx1078, nx1082, nx1084, nx1100, nx1110, nx1128, nx1130, nx1134, 
      nx1138, nx1140, nx1148, nx1154, nx1158, nx1174, nx1176, nx1186, nx1188, 
      nx1192, nx1202, nx1206, nx1216, nx1220, nx1230, nx1234, nx1244, nx1248, 
      nx1258, nx1262, nx1272, nx1276, nx1286, nx1290, nx1300, nx1304, nx1314, 
      nx1318, nx1328, nx1332, nx1342, nx1346, nx1356, nx1360, nx1370, nx1374, 
      nx1386, nx1388, nx1394, nx1398, nx1410, nx1422, nx1434, nx1446, nx1458, 
      nx1470, nx1482, nx1494, nx1506, nx1518, nx1530, nx1542, nx1554, 
      i5_MARo_0, i5_FAEN, nx1566, nx1576, nx1598, nx1604, nx1606, nx1614, 
      nx1616, nx1626, nx1634, nx1642, i5_MARo_1, nx1660, nx1668, nx1670, 
      i5_MARo_2, nx1682, nx1688, nx1696, nx1698, i5_MARo_3, nx1708, nx1716, 
      nx1724, nx1726, i5_MARo_4, nx1736, nx1744, nx1752, nx1754, i5_MARo_5, 
      nx1764, nx1772, nx1780, nx1782, i5_MARo_6, nx1794, nx1800, nx1808, 
      nx1810, i5_MARo_7, nx1820, nx1828, nx1836, nx1838, i5_MARo_8, nx1848, 
      nx1856, nx1864, nx1866, i5_MARo_9, nx1876, nx1884, nx1892, nx1894, 
      i5_MARo_10, nx1906, nx1912, nx1920, nx1922, i5_MARo_11, nx1932, nx1940, 
      nx1948, nx1950, i5_MARo_12, nx1960, nx1968, nx1976, nx1978, i5_MARo_13, 
      nx1988, nx1996, nx2004, nx2006, i5_MARo_14, nx2018, nx2024, nx2032, 
      nx2034, i5_MARo_15, nx2044, nx2052, nx2060, nx2062, nx2068, nx2072, 
      nx2080, nx2086, nx2098, nx2106, nx2108, nx2118, nx2122, nx2134, nx2148, 
      nx2160, nx2174, nx2186, nx2200, nx2212, nx2226, nx2238, nx2252, nx2264, 
      nx2278, nx2290, nx2304, nx2320, nx2334, nx2358, nx2382, nx2406, nx2430, 
      nx2444, nx2494, nx2512, nx2514, nx2520, nx2524, nx2548, nx2572, nx2596, 
      nx2620, nx2644, nx2668, nx2692, nx2708, nx2722, nx2746, nx2770, nx2794, 
      nx2818, nx2832, nx2880, nx2888, nx2902, nx2904, nx2910, nx2914, nx2938, 
      nx2962, nx2986, nx3010, nx3034, nx3058, nx3082, nx3098, nx3112, nx3136, 
      nx3160, nx3184, nx3208, nx3222, nx3272, nx3290, nx3292, nx3298, nx3302, 
      nx3326, nx3350, nx3374, nx3398, nx3422, nx3446, nx3470, nx3486, nx3500, 
      nx3524, nx3548, nx3572, nx3596, nx3610, nx3660, nx3668, nx3682, nx3686, 
      nx3688, nx3698, nx3702, nx3726, nx3750, nx3774, nx3798, nx3822, nx3846, 
      nx3870, nx3886, nx3900, nx3924, nx3948, nx3972, nx3996, nx4010, nx4060, 
      nx4074, nx4076, nx4082, nx4086, nx4110, nx4134, nx4158, nx4182, nx4206, 
      nx4230, nx4254, nx4270, nx4284, nx4308, nx4332, nx4356, nx4380, nx4394, 
      nx4446, nx4454, nx4468, nx4470, nx4476, nx4480, nx4504, nx4528, nx4552, 
      nx4576, nx4600, nx4624, nx4648, nx4664, nx4678, nx4702, nx4726, nx4750, 
      nx4774, nx4788, nx4838, nx4852, nx4854, nx4860, nx4864, nx4888, nx4912, 
      nx4936, nx4960, nx4984, nx5008, nx5032, nx5048, nx5062, nx5086, nx5110, 
      nx5134, nx5158, nx5172, nx5220, nx5228, nx5242, nx5246, nx5248, nx5258, 
      nx5262, nx5286, nx5310, nx5334, nx5358, nx5382, nx5406, nx5430, nx5446, 
      nx5460, nx5484, nx5508, nx5532, nx5556, nx5570, nx5620, nx5634, nx5636, 
      nx5642, nx5646, nx5670, nx5694, nx5718, nx5742, nx5766, nx5790, nx5814, 
      nx5830, nx5844, nx5868, nx5892, nx5916, nx5940, nx5954, nx6002, nx6010, 
      nx6024, nx6026, nx6032, nx6036, nx6060, nx6084, nx6108, nx6132, nx6156, 
      nx6180, nx6204, nx6220, nx6234, nx6258, nx6282, nx6306, nx6330, nx6344, 
      nx6394, nx6408, nx6410, nx6416, nx6420, nx6444, nx6468, nx6492, nx6516, 
      nx6540, nx6564, nx6588, nx6604, nx6618, nx6642, nx6666, nx6690, nx6714, 
      nx6728, nx6778, nx6786, nx6800, nx6802, nx6808, nx6812, nx6836, nx6860, 
      nx6884, nx6908, nx6932, nx6956, nx6980, nx6996, nx7010, nx7034, nx7058, 
      nx7082, nx7106, nx7120, nx7170, nx7184, nx7186, nx7192, nx7196, nx7220, 
      nx7244, nx7268, nx7292, nx7316, nx7340, nx7364, nx7380, nx7394, nx7418, 
      nx7442, nx7466, nx7490, nx7504, nx3127, nx3137, nx3147, nx3157, nx3167, 
      nx3177, nx3187, nx3197, nx3207, nx3217, nx3223, nx3225, nx3227, nx3233, 
      nx3235, nx3237, nx3247, nx3257, nx3267, nx3277, nx3283, nx3293, nx3307, 
      nx3317, nx3327, nx3337, nx3347, nx3357, nx3367, nx3377, nx3383, nx3393, 
      nx3407, nx3417, nx3427, nx3437, nx3447, nx3457, nx3467, nx3477, nx3483, 
      nx3493, nx3503, nx3518, nx3521, nx3523, nx3527, nx3533, nx3537, nx3541, 
      nx3545, nx3553, nx3555, nx3557, nx3561, nx3563, nx3565, nx3569, nx3571, 
      nx3575, nx3895, nx3899, nx3904, nx3907, nx3909, nx3917, nx3919, nx3921, 
      nx3925, nx3928, nx3930, nx3935, nx3938, nx3940, nx3943, nx3947, nx3955, 
      nx3959, nx3962, nx3967, nx3969, nx3971, nx3976, nx3979, nx3985, nx3988, 
      nx3993, nx3999, nx4002, nx4007, nx4011, nx4013, nx4016, nx4019, nx4022, 
      nx4026, nx4029, nx4033, nx4037, nx4041, nx4045, nx4050, nx4053, nx4059, 
      nx4063, nx4066, nx4073, nx4075, nx4079, nx4083, nx4090, nx4093, nx4100, 
      nx4107, nx4111, nx4114, nx4119, nx4124, nx4126, nx4131, nx4138, nx4141, 
      nx4148, nx4151, nx4155, nx4159, nx4162, nx4167, nx4171, nx4177, nx4179, 
      nx4181, nx4188, nx4191, nx4196, nx4198, nx4203, nx4207, nx4209, nx4212, 
      nx4215, nx4217, nx4220, nx4227, nx4231, nx4233, nx4237, nx4239, nx4243, 
      nx4246, nx4251, nx4255, nx4258, nx4261, nx4263, nx4267, nx4271, nx4274, 
      nx4277, nx4281, nx4283, nx4287, nx4293, nx4298, nx4301, nx4303, nx4307, 
      nx4309, nx4312, nx4315, nx4317, nx4318, nx4322, nx4327, nx4331, nx4333, 
      nx4336, nx4343, nx4345, nx4348, nx4353, nx4355, nx4359, nx4367, nx4370, 
      nx4374, nx4377, nx4379, nx4381, nx4383, nx4386, nx4389, nx4393, nx4397, 
      nx4399, nx4403, nx4405, nx4407, nx4409, nx4413, nx4417, nx4419, nx4425, 
      nx4427, nx4430, nx4434, nx4437, nx4441, nx4445, nx4447, nx4453, nx4457, 
      nx4460, nx4462, nx4465, nx4469, nx4475, nx4479, nx4485, nx4487, nx4496, 
      nx4501, nx4509, nx4511, nx4517, nx4522, nx4525, nx4532, nx4535, nx4537, 
      nx4542, nx4547, nx4553, nx4558, nx4565, nx4570, nx4577, nx4582, nx4592, 
      nx4613, nx4615, nx4618, nx4621, nx4625, nx4663, nx4665, nx4668, nx4670, 
      nx4673, nx4711, nx4715, nx4717, nx4720, nx4757, nx4759, nx4763, nx4765, 
      nx4804, nx4807, nx4809, nx4847, nx4851, nx4853, nx4894, nx4897, nx4899, 
      nx4937, nx4939, nx4942, nx4945, nx4985, nx4988, nx4990, nx5029, nx5033, 
      nx5035, nx5075, nx5078, nx5080, nx5119, nx5121, nx5124, nx5126, nx5165, 
      nx5169, nx5171, nx5209, nx5212, nx5215, nx5259, nx5263, nx5266, nx5303, 
      nx5305, nx5331, nx5333, nx5347, nx5349, nx5362, nx5375, nx5389, nx5403, 
      nx5415, nx5427, nx5441, nx5454, nx5467, nx5481, nx5497, nx5509, nx5522, 
      nx5535, nx5549, nx5562, nx5576, nx5589, nx5603, nx5615, nx5628, nx5643, 
      nx5659, nx5671, nx5684, nx5695, nx5697, nx5700, nx5703, nx5707, nx5709, 
      nx5712, nx5715, nx5719, nx5721, nx5724, nx5727, nx5731, nx5733, nx5736, 
      nx5739, nx5743, nx5745, nx5748, nx5751, nx5755, nx5757, nx5760, nx5763, 
      nx5767, nx5769, nx5772, nx5775, nx5779, nx5782, nx5785, nx5787, nx5791, 
      nx5793, nx5796, nx5799, nx5803, nx5805, nx5808, nx5811, nx5815, nx5817, 
      nx5820, nx5823, nx5827, nx5829, nx5833, nx5835, nx5838, nx5841, nx5845, 
      nx5847, nx5850, nx5853, nx5857, nx5859, nx5862, nx5865, nx5869, nx5872, 
      nx5875, nx5877, nx5881, nx5883, nx5886, nx5889, nx5893, nx5895, nx5898, 
      nx5901, nx5905, nx5907, nx5910, nx5913, nx5917, nx5919, nx5922, nx5925, 
      nx5929, nx5931, nx5934, nx5937, nx5941, nx5943, nx5946, nx5949, nx5953, 
      nx5955, nx5958, nx5961, nx5965, nx5967, nx5970, nx5973, nx5977, nx5979, 
      nx5982, nx5985, nx5989, nx5991, nx5994, nx5997, nx6001, nx6003, nx6007, 
      nx6009, nx6013, nx6015, nx6018, nx6021, nx6025, nx6027, nx6031, nx6033, 
      nx6037, nx6039, nx6042, nx6045, nx6049, nx6052, nx6055, nx6057, nx6061, 
      nx6063, nx6066, nx6069, nx6073, nx6075, nx6078, nx6081, nx6085, nx6087, 
      nx6090, nx6093, nx6097, nx6099, nx6102, nx6105, nx6109, nx6111, nx6114, 
      nx6117, nx6121, nx6123, nx6126, nx6129, nx6133, nx6135, nx6138, nx6141, 
      nx6145, nx6147, nx6150, nx6153, nx6157, nx6159, nx6162, nx6165, nx6169, 
      nx6171, nx6174, nx6177, nx6181, nx6183, nx6186, nx6189, nx6193, nx6195, 
      nx6198, nx6201, nx6205, nx6207, nx6210, nx6213, nx6217, nx6219, nx6223, 
      nx6225, nx6228, nx6231, nx6235, nx6237, nx6240, nx6243, nx6247, nx6249, 
      nx6252, nx6255, nx6259, nx6261, nx6264, nx6267, nx6271, nx6273, nx6276, 
      nx6279, nx6283, nx6285, nx6288, nx6291, nx6295, nx6297, nx6300, nx6303, 
      nx6307, nx6309, nx6312, nx6315, nx6319, nx6322, nx6325, nx6327, nx6331, 
      nx6333, nx6336, nx6339, nx6343, nx6345, nx6348, nx6350, nx6353, nx6355, 
      nx6358, nx6360, nx6363, nx6365, nx6368, nx6370, nx6373, nx6375, nx6379, 
      nx6381, nx6384, nx6387, nx6391, nx6393, nx6397, nx6399, nx6402, nx6405, 
      nx6409, nx6411, nx6415, nx6417, nx6421, nx6423, nx6426, nx6429, nx6433, 
      nx6435, nx6438, nx6441, nx6445, nx6447, nx6450, nx6453, nx6457, nx6459, 
      nx6462, nx6465, nx6469, nx6471, nx6474, nx6477, nx6481, nx6483, nx6486, 
      nx6489, nx6493, nx6496, nx6499, nx6501, nx6505, nx6507, nx6510, nx6513, 
      nx6517, nx6519, nx6522, nx6525, nx6529, nx6531, nx6534, nx6537, nx6541, 
      nx6543, nx6546, nx6549, nx6553, nx6555, nx6558, nx6561, nx6565, nx6567, 
      nx6570, nx6573, nx6577, nx6579, nx6582, nx6585, nx6589, nx6591, nx6594, 
      nx6597, nx6601, nx6603, nx6607, nx6609, nx6612, nx6615, nx6619, nx6621, 
      nx6624, nx6627, nx6631, nx6633, nx6636, nx6639, nx6643, nx6645, nx6648, 
      nx6651, nx6655, nx6657, nx6660, nx6663, nx6667, nx6669, nx6672, nx6675, 
      nx6679, nx6681, nx6684, nx6687, nx6691, nx6693, nx6696, nx6699, nx6703, 
      nx6705, nx6708, nx6711, nx6715, nx6717, nx6720, nx6723, nx6727, nx6729, 
      nx6732, nx6734, nx6737, nx6739, nx6742, nx6744, nx6747, nx6749, nx6752, 
      nx6754, nx6757, nx6761, nx6764, nx6766, nx6769, nx6771, nx6775, nx6777, 
      nx6781, nx6783, nx6787, nx6789, nx6792, nx6794, nx6797, nx6799, nx6803, 
      nx6805, nx6809, nx6811, nx6815, nx6817, nx6821, nx6823, nx6826, nx6828, 
      nx6831, nx6833, nx6837, nx6839, nx6842, nx6845, nx6849, nx6851, nx6854, 
      nx6857, nx6861, nx6863, nx6866, nx6869, nx6873, nx6875, nx6878, nx6881, 
      nx6885, nx6887, nx6890, nx6893, nx6897, nx6899, nx6902, nx6905, nx6909, 
      nx6911, nx6914, nx6917, nx6921, nx6923, nx6926, nx6929, nx6933, nx6936, 
      nx6939, nx6943, nx6946, nx6949, nx6953, nx6957, nx6960, nx6963, nx6967, 
      nx6970, nx6973, nx6977, nx6981, nx6984, nx6987, nx6991, nx6995, nx6999, 
      nx7002, nx7005, nx7009, nx7013, nx7016, nx7019, nx7023, nx7026, nx7029, 
      nx7033, nx7037, nx7039, nx7045, nx7048, nx7051, nx7057, nx7063, nx7067, 
      nx7072, nx7079, nx7081, nx7085, nx7088, nx7095, nx7098, nx7100, nx7103, 
      nx7107, nx7109, nx7115, nx7117, nx7121, nx7123, nx7126, nx7129, nx7132, 
      nx7137, nx7139, nx7143, nx7145, nx7148, nx7151, nx7157, nx7159, nx7163, 
      nx7165, nx7169, nx7173, nx7178, nx7181, nx7185, nx7189, nx7197, nx7199, 
      nx7202, nx7205, nx7209, nx7211, nx7214, nx7221, nx7223, nx7226, nx7229, 
      nx7233, nx7236, nx7241, nx7243, nx7247, nx7249, nx7253, nx7257, nx7262, 
      nx7265, nx7269, nx7272, nx7277, nx7279, nx7282, nx7284, nx7287, nx7289, 
      nx7293, nx7298, nx7301, nx7305, nx7307, nx7310, nx7313, nx7319, nx7321, 
      nx7325, nx7327, nx7330, nx7333, nx7339, nx7341, nx7344, nx7347, nx7354, 
      nx7356, nx7359, nx7361, nx7365, nx7367, nx7370, nx7377, nx7381, nx7383, 
      nx7390, nx7392, nx7395, nx7397, nx7399, nx7401, nx7403, nx7405, nx7407, 
      nx7409, nx7411, nx7413, nx7415, nx7417, nx7419, nx7421, nx7423, nx7425, 
      nx7427, nx7429, nx7431, nx7433, nx7435, nx7437, nx7439, nx7441, nx7443, 
      nx7445, nx7447, nx7449, nx7451, nx7455, nx7457, nx7459, nx7461, nx7463, 
      nx7465, nx7467, nx7469, nx7471, nx7473, nx7475, nx7477, nx7479, nx7481, 
      nx7483, nx7485, nx7487, nx7489, nx7491, nx7493, nx7495, nx7497, nx7499, 
      nx7501, nx7503, nx7505, nx7507, nx7509, nx7511, nx7515, nx7517, nx7519, 
      nx7521, nx7523, nx7525, nx7527, nx7529, nx7531, nx7537, nx7539, nx7541, 
      nx7551, nx7553, nx7555, nx7557, nx7559, nx7561, nx7563, nx7565, nx7567, 
      nx7569, nx7571, nx7575, nx7577, nx7579, nx7581, nx7583, nx7587, nx7589, 
      nx7591, nx7593, nx7595, nx7599, nx7601, nx7603, nx7605, nx7607, nx7611, 
      nx7613, nx7615, nx7617, nx7619, nx7623, nx7625, nx7627, nx7629, nx7631, 
      nx7633, nx7635, nx7637, nx7639, nx7643, nx7645, nx7647, nx7649, nx7651, 
      nx7655, nx7657, nx7659, nx7661, nx7663, nx7667, nx7669, nx7671, nx7673, 
      nx7675, nx7679, nx7681, nx7683, nx7685, nx7687, nx7691, nx7693, nx7695, 
      nx7697, nx7699, nx7703, nx7705, nx7707, nx7709, nx7711, nx7715, nx7717, 
      nx7719, nx7721, nx7723, nx7727, nx7729, nx7731, nx7733, nx7735, nx7737, 
      nx7739, nx7741, nx7743, nx7745, nx7747, nx7749, nx7751, nx7753, nx7755, 
      nx7757, nx7759, nx7761, nx7763, nx7765, nx7767, nx7769, nx7771, nx7773, 
      nx7775, nx7777, nx7779, nx7781, nx7783, nx7785, nx7787, nx7789, nx7791, 
      nx7793, nx7795, nx7797, nx7799, nx7801, nx7803, nx7805, nx7807, nx7809, 
      nx7811, nx7813, nx7815, nx7817, nx7819, nx7821, nx7823, nx7825, nx7827, 
      nx7829, nx7831, nx7833, nx7835, nx7837, nx7839, nx7841, nx7843, nx7845, 
      nx7847, nx7849, nx7851, nx7853, nx7855, nx7857, nx7859, nx7861, nx7863, 
      nx7865, nx7867, nx7869, nx7871, nx7873, nx7875, nx7877, nx7879, nx7881, 
      nx7883, nx7885, nx7887, nx7889, nx7891, nx7893, nx7895, nx7897, nx7899, 
      nx7901, nx7907, nx7909, nx7911, nx7913, nx7957, nx7959, nx7961, nx8009, 
      nx8011, nx8013, nx8015, nx8017, nx8019, nx8021, nx8023, nx8025, nx8027, 
      nx8029, nx8031, nx8033, nx8035, nx8037, nx8039, nx8041, nx8043, nx8045, 
      nx8047, nx8049, nx8051, nx8053, nx8055, nx8057, nx8059, nx8061, nx8063, 
      nx8065, nx8067, nx8069, nx8071, nx8073, nx8075, nx8077, nx8079, nx8081, 
      nx8083, nx8085, nx8087, nx8089, nx5, nx8093, nx8096, nx8099, nx8102, 
      nx8105, nx8108, nx8111, nx8114, nx8117, nx8120, nx8123, nx8126, nx8129, 
      nx8132, nx8135, nx8138, nx8141, nx8144, nx8147, nx8150, nx8153, nx8156, 
      nx8159, nx8162, nx8165, nx8168, nx8171, nx8174, nx8177, nx8180, nx8183, 
      nx8186, nx8189, nx8192, nx8195, nx8198, nx8201, nx8204, nx8207, nx8210, 
      nx8213, nx8216, nx8219, nx8222, nx8225, nx8228, nx8231, nx8234, nx8237, 
      nx8240, nx8243, nx8246, nx8249, nx8252, nx8255, nx8258, nx8261, nx8264, 
      nx8267, nx8270, nx8273, nx8276, nx8279, nx8282, nx8285, nx8288, nx8291, 
      nx8294, nx8297, nx8300, nx8303, nx8306, nx8309, nx8312, nx8315, nx8318, 
      nx8321, nx8324, nx8327, nx8330, nx8333, nx8336, nx8339, nx8342, nx8345, 
      nx8348, nx8351, nx8354, nx8357, nx8360, nx8363, nx8366, nx8369, nx8372, 
      nx8375, nx8378, nx8381, nx8384, nx8387, nx8390, nx8393, nx8396, nx8399, 
      nx8402, nx8405, nx8408, nx8411, nx8414, nx8417, nx8420, nx8423, nx8426, 
      nx8429, nx8432, nx8435, nx8438, nx8441, nx8444, nx8447, nx8450, nx8453, 
      nx8456, nx8459, nx8462, nx8465, nx8468, nx8471, nx8474, nx8477, nx8480, 
      nx8483, nx8486, nx8489, nx8492, nx8495, nx8498, nx8501, nx8504, nx8507, 
      nx8510, nx8513, nx8516, nx8519, nx8522, nx8525, nx8528, nx8531, nx8534, 
      nx8537, nx8540, nx8543, nx8546, nx8549, nx8552, nx8555, nx8558, nx8561, 
      nx8564, nx8567, nx8570, nx8573, nx8576, nx8579, nx8582, nx8585, nx8588, 
      nx8591, nx8594, nx8597, nx8600, nx8603, nx8606, nx8609, nx8612, nx8615, 
      nx8618, nx8621, nx8624, nx8627, nx8630, nx8633, nx8636, nx8639, nx8642, 
      nx8645, nx8648, nx8651, nx8654, nx8657, nx8660, nx8663, nx8666, nx8669, 
      nx8672, nx8675, nx8678, nx8681, nx8684, nx8687, nx8690, nx8693, nx8696, 
      nx8699, nx8702, nx8705, nx8708, nx8711, nx8714, nx8717, nx8720, nx8723, 
      nx8726, nx8729, nx8732, nx8735, nx8738, nx8741, nx8744, nx8747, nx8750, 
      nx8753, nx8756, nx8759, nx8762, nx8765, nx8768, nx8771, nx8774, nx8777, 
      nx8780, nx8783, nx8786, nx8789, nx8792, nx8795, nx8798, nx8801, nx8804, 
      nx8807, nx8810, nx8813, nx8816, nx8819, nx8822, nx8825, nx8828, nx8831, 
      nx8834, nx8837, nx8840, nx8843, nx8846, nx8849, nx8852, nx8855, nx8858, 
      nx8861, nx8864, nx8867, nx8870, nx8873, nx8876, nx8879, nx8882, nx8885, 
      nx8888, nx8891, nx8894, nx8897, nx8900, nx8903, nx8906, nx8909, nx8912, 
      nx8915, nx8918, nx8921, nx8924, nx8927, nx8930, nx8933, nx8936, nx8939, 
      nx8942, nx8945, nx8948, nx8951, nx8954, nx8957, nx8960, nx8963, nx8966, 
      nx8969, nx8972, nx8975, nx8978, nx8981, nx8984, nx8987, nx8990, nx8993, 
      nx8996, nx8999, nx9002, nx9005, nx9008, nx9011, nx9014, nx9017, nx9020, 
      nx9023, nx9026, nx9029, nx9032, nx9035, nx9038, nx9041, nx9044, nx9047, 
      nx9050, nx9053, nx9056, nx9059, nx9062, nx9065, nx9068, nx9071, nx9074, 
      nx9077, nx9080, nx9083, nx9086, nx9089, nx9092, nx9095, nx9098, nx9101, 
      nx9104, nx9107, nx9110, nx9113, nx9116, nx9119, nx9122, nx9125, nx9128, 
      nx9131, nx9134, nx9137, nx9140, nx9143, nx9146, nx9149, nx9152, nx9155, 
      nx9158, nx9161, nx9164, nx9167, nx9170, nx9173, nx9176, nx9179, nx9182, 
      nx9185, nx9188, nx9191, nx9194, nx9197, nx9200, nx9203, nx9206, nx9209, 
      nx9212, nx9215, nx9218, nx9221, nx9224, nx9227, nx9230, nx9233, nx9236, 
      nx9239, nx9242, nx9245, nx9248, nx9251, nx9254, nx9257, nx9260, nx9263, 
      nx9266, nx9269, nx9272, nx9274, nx9276, nx9278, nx9280, nx9282, nx9284, 
      nx9286, nx9288, nx9290, nx9292, nx9294, nx9296, nx9298, nx9300, nx9302, 
      nx9304, nx9306, nx9308, nx9310, nx9312, nx9314, nx9316, nx9318, nx9320, 
      nx9322, nx9324, nx9326, nx9328, nx9330, nx9332, nx9334, nx9336, nx9338, 
      nx9340, nx9342, nx9344, nx9346, nx9348, nx9350, nx9352, nx9354, nx9356, 
      nx9358, nx9360, nx9362, nx9364, nx9366, nx9368, nx9370, nx9372, nx9374, 
      nx9376, nx9378, nx9380, nx9382, nx9384, nx9386, nx9388, nx9390, nx9392, 
      nx9394, nx9396, nx9398, nx9400, nx9402, nx9404, nx9406, nx9408: 
   std_logic ;

begin
   Result(3) <= ResultIn(3) ;
   Result(2) <= ResultIn(2) ;
   Result(1) <= ResultIn(1) ;
   Result(0) <= ResultIn(0) ;
   DecompressedData(254) <= DecompressedData(255) ;
   DecompressedData(253) <= DecompressedData(255) ;
   DecompressedData(238) <= DecompressedData(239) ;
   DecompressedData(237) <= DecompressedData(239) ;
   DecompressedData1(254) <= DecompressedData1(255) ;
   DecompressedData1(253) <= DecompressedData1(255) ;
   DecompressedData1(252) <= DecompressedData1(255) ;
   DecompressedData1(251) <= DecompressedData1(255) ;
   DecompressedData1(250) <= DecompressedData1(255) ;
   DecompressedData1(249) <= DecompressedData1(255) ;
   DecompressedData1(248) <= DecompressedData1(255) ;
   DecompressedData1(247) <= DecompressedData1(255) ;
   DecompressedData1(246) <= DecompressedData1(255) ;
   DecompressedData1(245) <= DecompressedData1(255) ;
   DecompressedData1(244) <= DecompressedData1(255) ;
   DecompressedData1(243) <= DecompressedData1(255) ;
   DecompressedData1(242) <= DecompressedData1(255) ;
   DecompressedData1(241) <= DecompressedData1(255) ;
   DecompressedData1(240) <= DecompressedData1(255) ;
   DecompressedData1(239) <= DecompressedData1(255) ;
   DecompressedData1(238) <= DecompressedData1(255) ;
   DecompressedData1(237) <= DecompressedData1(255) ;
   DecompressedData1(236) <= DecompressedData1(255) ;
   DecompressedData1(235) <= DecompressedData1(255) ;
   DecompressedData1(234) <= DecompressedData1(255) ;
   DecompressedData1(233) <= DecompressedData1(255) ;
   DecompressedData1(232) <= DecompressedData1(255) ;
   DecompressedData1(231) <= DecompressedData1(255) ;
   DecompressedData1(230) <= DecompressedData1(255) ;
   DecompressedData1(229) <= DecompressedData1(255) ;
   DecompressedData1(228) <= DecompressedData1(255) ;
   DecompressedData1(227) <= DecompressedData1(255) ;
   DecompressedData1(226) <= DecompressedData1(255) ;
   DecompressedData1(225) <= DecompressedData1(255) ;
   DecompressedData1(224) <= DecompressedData1(255) ;
   DecompressedData2(254) <= DecompressedData2(255) ;
   DecompressedData2(253) <= DecompressedData2(255) ;
   DecompressedData2(238) <= DecompressedData2(239) ;
   DecompressedData2(237) <= DecompressedData2(239) ;
   DecompressedData2(222) <= DecompressedData2(223) ;
   DecompressedData2(221) <= DecompressedData2(223) ;
   DecompressedData2(206) <= DecompressedData2(207) ;
   DecompressedData2(205) <= DecompressedData2(207) ;
   DecompressedData2(190) <= DecompressedData2(191) ;
   DecompressedData2(189) <= DecompressedData2(191) ;
   DecompressedData2(174) <= DecompressedData2(175) ;
   DecompressedData2(173) <= DecompressedData2(175) ;
   DecompressedData2(158) <= DecompressedData2(159) ;
   DecompressedData2(157) <= DecompressedData2(159) ;
   DecompressedData2(142) <= DecompressedData2(143) ;
   DecompressedData2(141) <= DecompressedData2(143) ;
   DecompressedData2(126) <= DecompressedData2(127) ;
   DecompressedData2(125) <= DecompressedData2(127) ;
   DecompressedData2(110) <= DecompressedData2(111) ;
   DecompressedData2(109) <= DecompressedData2(111) ;
   DecompressedData2(94) <= DecompressedData2(95) ;
   DecompressedData2(93) <= DecompressedData2(95) ;
   DecompressedData2(78) <= DecompressedData2(79) ;
   DecompressedData2(77) <= DecompressedData2(79) ;
   DecompressedData2(62) <= DecompressedData2(63) ;
   DecompressedData2(61) <= DecompressedData2(63) ;
   DecompressedData2(46) <= DecompressedData2(47) ;
   DecompressedData2(45) <= DecompressedData2(47) ;
   DecompressedData2(30) <= DecompressedData2(31) ;
   DecompressedData2(29) <= DecompressedData2(31) ;
   DecompressedData2(14) <= DecompressedData2(15) ;
   DecompressedData2(13) <= DecompressedData2(15) ;
   PClk <= CLK ;
   ProcessEnable <= ProcessEnable_EXMPLR ;
   ix3 : fake_vcc port map ( Y=>nx2);
   ix2589 : fake_gnd port map ( Y=>DecompressedData1(255));
   ix631 : nor02_2x port map ( Y=>loadingimg, A0=>CNNIMGLOAD, A1=>nx7957);
   ix83 : nor02_2x port map ( Y=>nx82, A0=>LP, A1=>nx3518);
   ix3519 : nor02_2x port map ( Y=>nx3518, A0=>nx74, A1=>nx7737);
   ix75 : nor02_2x port map ( Y=>nx74, A0=>nx3521, A1=>Rst);
   ix3522 : inv01 port map ( Y=>nx3521, A=>INTR);
   ix67 : nor02_2x port map ( Y=>nx66, A0=>nx3527, A1=>nx3533);
   ix3528 : nand04 port map ( Y=>nx3527, A0=>nx8, A1=>nx14, A2=>nx22, A3=>
      nx28);
   ix9 : nor02_2x port map ( Y=>nx8, A0=>DataBus(8), A1=>DataBus(9));
   ix15 : nor02_2x port map ( Y=>nx14, A0=>DataBus(10), A1=>DataBus(11));
   ix23 : nor02_2x port map ( Y=>nx22, A0=>DataBus(12), A1=>DataBus(13));
   ix29 : nor02_2x port map ( Y=>nx28, A0=>DataBus(0), A1=>DataBus(1));
   ix3534 : nand04 port map ( Y=>nx3533, A0=>nx46, A1=>nx52, A2=>nx3541, A3
      =>nx7907);
   ix47 : nor03_2x port map ( Y=>nx46, A0=>DataBus(2), A1=>DataBus(3), A2=>
      nx3537);
   ix3538 : inv01 port map ( Y=>nx3537, A=>nx44);
   ix45 : nor02_2x port map ( Y=>nx44, A0=>DataBus(4), A1=>DataBus(5));
   ix53 : nor02_2x port map ( Y=>nx52, A0=>DataBus(6), A1=>DataBus(7));
   ix3542 : nor02_2x port map ( Y=>nx3541, A0=>DataBus(14), A1=>DataBus(15)
   );
   i1_L_reg_Q : dff port map ( Q=>loadenable, QB=>OPEN, D=>nx82, CLK=>nx70);
   ix71 : nand02 port map ( Y=>nx70, A0=>nx7737, A1=>nx3521);
   ix3546 : inv01 port map ( Y=>nx3545, A=>Rst);
   ix91 : nor02_2x port map ( Y=>loadingCNN, A0=>nx7741, A1=>nx7957);
   i0_L_reg_Q : dff port map ( Q=>ProcessEnable_EXMPLR, QB=>nx3563, D=>
      nx1576, CLK=>nx1566);
   ix1577 : nor02_2x port map ( Y=>nx1576, A0=>nx3553, A1=>nx3557);
   ix3554 : nor02_2x port map ( Y=>nx3553, A0=>nx3555, A1=>INTR);
   ix3556 : inv01 port map ( Y=>nx3555, A=>PDone);
   ix3558 : nand02 port map ( Y=>nx3557, A0=>LP, A1=>nx3545);
   ix1567 : nand02 port map ( Y=>nx1566, A0=>nx3561, A1=>nx3545);
   ix3562 : nor02_2x port map ( Y=>nx3561, A0=>PDone, A1=>INTR);
   ix7553 : nand02 port map ( Y=>Done, A0=>nx3565, A1=>nx3555);
   ix3566 : nand03 port map ( Y=>nx3565, A0=>nx32, A1=>nx46, A2=>nx62);
   ix33 : nor02_2x port map ( Y=>nx32, A0=>nx3569, A1=>nx3571);
   ix3570 : nand02 port map ( Y=>nx3569, A0=>nx8, A1=>nx14);
   ix3572 : nand02 port map ( Y=>nx3571, A0=>nx22, A1=>nx28);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>DataBus(6), A1=>DataBus(7), A2=>
      nx3575);
   ix3576 : nand02 port map ( Y=>nx3575, A0=>nx3541, A1=>nx7907);
   tri_DataFromRam_0 : tri01 port map ( Y=>DataFromRam(0), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_1 : tri01 port map ( Y=>DataFromRam(1), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_2 : tri01 port map ( Y=>DataFromRam(2), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_3 : tri01 port map ( Y=>DataFromRam(3), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_4 : tri01 port map ( Y=>DataFromRam(4), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_5 : tri01 port map ( Y=>DataFromRam(5), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_6 : tri01 port map ( Y=>DataFromRam(6), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_7 : tri01 port map ( Y=>DataFromRam(7), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_8 : tri01 port map ( Y=>DataFromRam(8), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_9 : tri01 port map ( Y=>DataFromRam(9), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_10 : tri01 port map ( Y=>DataFromRam(10), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_11 : tri01 port map ( Y=>DataFromRam(11), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_12 : tri01 port map ( Y=>DataFromRam(12), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_13 : tri01 port map ( Y=>DataFromRam(13), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_14 : tri01 port map ( Y=>DataFromRam(14), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_15 : tri01 port map ( Y=>DataFromRam(15), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_16 : tri01 port map ( Y=>DataFromRam(16), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_17 : tri01 port map ( Y=>DataFromRam(17), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_18 : tri01 port map ( Y=>DataFromRam(18), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_19 : tri01 port map ( Y=>DataFromRam(19), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_20 : tri01 port map ( Y=>DataFromRam(20), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_21 : tri01 port map ( Y=>DataFromRam(21), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_22 : tri01 port map ( Y=>DataFromRam(22), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_23 : tri01 port map ( Y=>DataFromRam(23), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_24 : tri01 port map ( Y=>DataFromRam(24), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_25 : tri01 port map ( Y=>DataFromRam(25), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_26 : tri01 port map ( Y=>DataFromRam(26), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_27 : tri01 port map ( Y=>DataFromRam(27), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_28 : tri01 port map ( Y=>DataFromRam(28), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_29 : tri01 port map ( Y=>DataFromRam(29), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_30 : tri01 port map ( Y=>DataFromRam(30), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_31 : tri01 port map ( Y=>DataFromRam(31), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_32 : tri01 port map ( Y=>DataFromRam(32), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_33 : tri01 port map ( Y=>DataFromRam(33), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_34 : tri01 port map ( Y=>DataFromRam(34), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_35 : tri01 port map ( Y=>DataFromRam(35), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_36 : tri01 port map ( Y=>DataFromRam(36), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_37 : tri01 port map ( Y=>DataFromRam(37), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_38 : tri01 port map ( Y=>DataFromRam(38), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_39 : tri01 port map ( Y=>DataFromRam(39), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_40 : tri01 port map ( Y=>DataFromRam(40), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_41 : tri01 port map ( Y=>DataFromRam(41), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_42 : tri01 port map ( Y=>DataFromRam(42), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_43 : tri01 port map ( Y=>DataFromRam(43), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_44 : tri01 port map ( Y=>DataFromRam(44), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_45 : tri01 port map ( Y=>DataFromRam(45), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_46 : tri01 port map ( Y=>DataFromRam(46), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_47 : tri01 port map ( Y=>DataFromRam(47), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_48 : tri01 port map ( Y=>DataFromRam(48), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_49 : tri01 port map ( Y=>DataFromRam(49), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_50 : tri01 port map ( Y=>DataFromRam(50), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_51 : tri01 port map ( Y=>DataFromRam(51), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_52 : tri01 port map ( Y=>DataFromRam(52), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_53 : tri01 port map ( Y=>DataFromRam(53), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_54 : tri01 port map ( Y=>DataFromRam(54), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_55 : tri01 port map ( Y=>DataFromRam(55), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_56 : tri01 port map ( Y=>DataFromRam(56), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_57 : tri01 port map ( Y=>DataFromRam(57), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_58 : tri01 port map ( Y=>DataFromRam(58), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_59 : tri01 port map ( Y=>DataFromRam(59), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_60 : tri01 port map ( Y=>DataFromRam(60), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_61 : tri01 port map ( Y=>DataFromRam(61), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_62 : tri01 port map ( Y=>DataFromRam(62), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_63 : tri01 port map ( Y=>DataFromRam(63), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_64 : tri01 port map ( Y=>DataFromRam(64), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_65 : tri01 port map ( Y=>DataFromRam(65), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_66 : tri01 port map ( Y=>DataFromRam(66), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_67 : tri01 port map ( Y=>DataFromRam(67), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_68 : tri01 port map ( Y=>DataFromRam(68), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_69 : tri01 port map ( Y=>DataFromRam(69), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_70 : tri01 port map ( Y=>DataFromRam(70), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_71 : tri01 port map ( Y=>DataFromRam(71), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_72 : tri01 port map ( Y=>DataFromRam(72), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_73 : tri01 port map ( Y=>DataFromRam(73), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_74 : tri01 port map ( Y=>DataFromRam(74), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_75 : tri01 port map ( Y=>DataFromRam(75), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_76 : tri01 port map ( Y=>DataFromRam(76), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_77 : tri01 port map ( Y=>DataFromRam(77), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_78 : tri01 port map ( Y=>DataFromRam(78), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_79 : tri01 port map ( Y=>DataFromRam(79), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_80 : tri01 port map ( Y=>DataFromRam(80), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_81 : tri01 port map ( Y=>DataFromRam(81), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_82 : tri01 port map ( Y=>DataFromRam(82), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_83 : tri01 port map ( Y=>DataFromRam(83), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_84 : tri01 port map ( Y=>DataFromRam(84), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_85 : tri01 port map ( Y=>DataFromRam(85), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_86 : tri01 port map ( Y=>DataFromRam(86), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_87 : tri01 port map ( Y=>DataFromRam(87), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_88 : tri01 port map ( Y=>DataFromRam(88), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_89 : tri01 port map ( Y=>DataFromRam(89), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_90 : tri01 port map ( Y=>DataFromRam(90), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_91 : tri01 port map ( Y=>DataFromRam(91), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_92 : tri01 port map ( Y=>DataFromRam(92), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_93 : tri01 port map ( Y=>DataFromRam(93), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_94 : tri01 port map ( Y=>DataFromRam(94), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_95 : tri01 port map ( Y=>DataFromRam(95), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_96 : tri01 port map ( Y=>DataFromRam(96), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_97 : tri01 port map ( Y=>DataFromRam(97), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_98 : tri01 port map ( Y=>DataFromRam(98), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_99 : tri01 port map ( Y=>DataFromRam(99), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_100 : tri01 port map ( Y=>DataFromRam(100), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_101 : tri01 port map ( Y=>DataFromRam(101), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_102 : tri01 port map ( Y=>DataFromRam(102), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_103 : tri01 port map ( Y=>DataFromRam(103), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_104 : tri01 port map ( Y=>DataFromRam(104), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_105 : tri01 port map ( Y=>DataFromRam(105), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_106 : tri01 port map ( Y=>DataFromRam(106), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_107 : tri01 port map ( Y=>DataFromRam(107), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_108 : tri01 port map ( Y=>DataFromRam(108), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_109 : tri01 port map ( Y=>DataFromRam(109), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_110 : tri01 port map ( Y=>DataFromRam(110), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_111 : tri01 port map ( Y=>DataFromRam(111), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_112 : tri01 port map ( Y=>DataFromRam(112), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_113 : tri01 port map ( Y=>DataFromRam(113), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_114 : tri01 port map ( Y=>DataFromRam(114), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_115 : tri01 port map ( Y=>DataFromRam(115), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_116 : tri01 port map ( Y=>DataFromRam(116), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_117 : tri01 port map ( Y=>DataFromRam(117), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_118 : tri01 port map ( Y=>DataFromRam(118), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_119 : tri01 port map ( Y=>DataFromRam(119), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_120 : tri01 port map ( Y=>DataFromRam(120), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_121 : tri01 port map ( Y=>DataFromRam(121), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_122 : tri01 port map ( Y=>DataFromRam(122), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_123 : tri01 port map ( Y=>DataFromRam(123), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_124 : tri01 port map ( Y=>DataFromRam(124), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_125 : tri01 port map ( Y=>DataFromRam(125), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_126 : tri01 port map ( Y=>DataFromRam(126), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_127 : tri01 port map ( Y=>DataFromRam(127), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_128 : tri01 port map ( Y=>DataFromRam(128), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_129 : tri01 port map ( Y=>DataFromRam(129), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_130 : tri01 port map ( Y=>DataFromRam(130), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_131 : tri01 port map ( Y=>DataFromRam(131), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_132 : tri01 port map ( Y=>DataFromRam(132), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_133 : tri01 port map ( Y=>DataFromRam(133), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_134 : tri01 port map ( Y=>DataFromRam(134), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_135 : tri01 port map ( Y=>DataFromRam(135), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_136 : tri01 port map ( Y=>DataFromRam(136), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_137 : tri01 port map ( Y=>DataFromRam(137), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_138 : tri01 port map ( Y=>DataFromRam(138), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_139 : tri01 port map ( Y=>DataFromRam(139), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_140 : tri01 port map ( Y=>DataFromRam(140), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_141 : tri01 port map ( Y=>DataFromRam(141), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_142 : tri01 port map ( Y=>DataFromRam(142), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_143 : tri01 port map ( Y=>DataFromRam(143), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_144 : tri01 port map ( Y=>DataFromRam(144), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_145 : tri01 port map ( Y=>DataFromRam(145), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_146 : tri01 port map ( Y=>DataFromRam(146), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_147 : tri01 port map ( Y=>DataFromRam(147), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_148 : tri01 port map ( Y=>DataFromRam(148), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_149 : tri01 port map ( Y=>DataFromRam(149), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_150 : tri01 port map ( Y=>DataFromRam(150), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_151 : tri01 port map ( Y=>DataFromRam(151), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_152 : tri01 port map ( Y=>DataFromRam(152), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_153 : tri01 port map ( Y=>DataFromRam(153), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_154 : tri01 port map ( Y=>DataFromRam(154), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_155 : tri01 port map ( Y=>DataFromRam(155), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_156 : tri01 port map ( Y=>DataFromRam(156), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_157 : tri01 port map ( Y=>DataFromRam(157), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_158 : tri01 port map ( Y=>DataFromRam(158), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_159 : tri01 port map ( Y=>DataFromRam(159), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_160 : tri01 port map ( Y=>DataFromRam(160), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_161 : tri01 port map ( Y=>DataFromRam(161), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_162 : tri01 port map ( Y=>DataFromRam(162), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_163 : tri01 port map ( Y=>DataFromRam(163), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_164 : tri01 port map ( Y=>DataFromRam(164), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_165 : tri01 port map ( Y=>DataFromRam(165), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_166 : tri01 port map ( Y=>DataFromRam(166), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_167 : tri01 port map ( Y=>DataFromRam(167), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_168 : tri01 port map ( Y=>DataFromRam(168), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_169 : tri01 port map ( Y=>DataFromRam(169), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_170 : tri01 port map ( Y=>DataFromRam(170), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_171 : tri01 port map ( Y=>DataFromRam(171), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_172 : tri01 port map ( Y=>DataFromRam(172), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_173 : tri01 port map ( Y=>DataFromRam(173), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_174 : tri01 port map ( Y=>DataFromRam(174), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_175 : tri01 port map ( Y=>DataFromRam(175), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_176 : tri01 port map ( Y=>DataFromRam(176), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_177 : tri01 port map ( Y=>DataFromRam(177), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_178 : tri01 port map ( Y=>DataFromRam(178), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_179 : tri01 port map ( Y=>DataFromRam(179), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_180 : tri01 port map ( Y=>DataFromRam(180), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_181 : tri01 port map ( Y=>DataFromRam(181), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_182 : tri01 port map ( Y=>DataFromRam(182), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_183 : tri01 port map ( Y=>DataFromRam(183), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_184 : tri01 port map ( Y=>DataFromRam(184), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_185 : tri01 port map ( Y=>DataFromRam(185), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_186 : tri01 port map ( Y=>DataFromRam(186), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_187 : tri01 port map ( Y=>DataFromRam(187), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_188 : tri01 port map ( Y=>DataFromRam(188), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_189 : tri01 port map ( Y=>DataFromRam(189), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_190 : tri01 port map ( Y=>DataFromRam(190), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_191 : tri01 port map ( Y=>DataFromRam(191), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_192 : tri01 port map ( Y=>DataFromRam(192), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_193 : tri01 port map ( Y=>DataFromRam(193), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_194 : tri01 port map ( Y=>DataFromRam(194), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_195 : tri01 port map ( Y=>DataFromRam(195), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_196 : tri01 port map ( Y=>DataFromRam(196), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_197 : tri01 port map ( Y=>DataFromRam(197), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_198 : tri01 port map ( Y=>DataFromRam(198), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_199 : tri01 port map ( Y=>DataFromRam(199), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_200 : tri01 port map ( Y=>DataFromRam(200), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_201 : tri01 port map ( Y=>DataFromRam(201), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_202 : tri01 port map ( Y=>DataFromRam(202), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_203 : tri01 port map ( Y=>DataFromRam(203), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_204 : tri01 port map ( Y=>DataFromRam(204), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_205 : tri01 port map ( Y=>DataFromRam(205), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_206 : tri01 port map ( Y=>DataFromRam(206), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_207 : tri01 port map ( Y=>DataFromRam(207), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_208 : tri01 port map ( Y=>DataFromRam(208), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_209 : tri01 port map ( Y=>DataFromRam(209), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_210 : tri01 port map ( Y=>DataFromRam(210), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_211 : tri01 port map ( Y=>DataFromRam(211), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_212 : tri01 port map ( Y=>DataFromRam(212), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_213 : tri01 port map ( Y=>DataFromRam(213), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_214 : tri01 port map ( Y=>DataFromRam(214), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_215 : tri01 port map ( Y=>DataFromRam(215), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_216 : tri01 port map ( Y=>DataFromRam(216), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_217 : tri01 port map ( Y=>DataFromRam(217), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_218 : tri01 port map ( Y=>DataFromRam(218), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_219 : tri01 port map ( Y=>DataFromRam(219), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_220 : tri01 port map ( Y=>DataFromRam(220), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_221 : tri01 port map ( Y=>DataFromRam(221), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_222 : tri01 port map ( Y=>DataFromRam(222), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_223 : tri01 port map ( Y=>DataFromRam(223), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_224 : tri01 port map ( Y=>DataFromRam(224), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_225 : tri01 port map ( Y=>DataFromRam(225), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_226 : tri01 port map ( Y=>DataFromRam(226), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_227 : tri01 port map ( Y=>DataFromRam(227), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_228 : tri01 port map ( Y=>DataFromRam(228), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_229 : tri01 port map ( Y=>DataFromRam(229), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_230 : tri01 port map ( Y=>DataFromRam(230), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_231 : tri01 port map ( Y=>DataFromRam(231), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_232 : tri01 port map ( Y=>DataFromRam(232), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_233 : tri01 port map ( Y=>DataFromRam(233), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_234 : tri01 port map ( Y=>DataFromRam(234), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_235 : tri01 port map ( Y=>DataFromRam(235), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_236 : tri01 port map ( Y=>DataFromRam(236), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_237 : tri01 port map ( Y=>DataFromRam(237), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_238 : tri01 port map ( Y=>DataFromRam(238), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_239 : tri01 port map ( Y=>DataFromRam(239), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_240 : tri01 port map ( Y=>DataFromRam(240), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_241 : tri01 port map ( Y=>DataFromRam(241), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_242 : tri01 port map ( Y=>DataFromRam(242), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_243 : tri01 port map ( Y=>DataFromRam(243), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_244 : tri01 port map ( Y=>DataFromRam(244), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_245 : tri01 port map ( Y=>DataFromRam(245), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_246 : tri01 port map ( Y=>DataFromRam(246), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_247 : tri01 port map ( Y=>DataFromRam(247), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_248 : tri01 port map ( Y=>DataFromRam(248), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_249 : tri01 port map ( Y=>DataFromRam(249), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_250 : tri01 port map ( Y=>DataFromRam(250), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_251 : tri01 port map ( Y=>DataFromRam(251), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_252 : tri01 port map ( Y=>DataFromRam(252), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_253 : tri01 port map ( Y=>DataFromRam(253), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_254 : tri01 port map ( Y=>DataFromRam(254), A=>nx2, E=>
      DecompressedData1(255));
   tri_DataFromRam_255 : tri01 port map ( Y=>DataFromRam(255), A=>nx2, E=>
      DecompressedData1(255));
   ix611 : aoi21 port map ( Y=>nx610, A0=>nx7765, A1=>zed, B0=>nx4198);
   ix3896 : nor02_2x port map ( Y=>nx3895, A0=>nx3093, A1=>nx282);
   ix191 : nand03 port map ( Y=>nx3093, A0=>nx3899, A1=>nx4019, A2=>nx4033);
   ix3900 : nor02_2x port map ( Y=>nx3899, A0=>i8_counterout1_0, A1=>
      i8_counterout1_1);
   ix3128 : oai21 port map ( Y=>nx3127, A0=>nx3904, A1=>nx7805, B0=>nx4196);
   ix3905 : nor02_2x port map ( Y=>nx3904, A0=>nx136, A1=>nx128);
   ix137 : oai21 port map ( Y=>nx136, A0=>nx3907, A1=>nx3909, B0=>nx4188);
   reg_i8_counterout1_0 : dff port map ( Q=>i8_counterout1_0, QB=>nx3907, D
      =>nx3127, CLK=>CLK);
   ix3910 : oai21 port map ( Y=>nx3909, A0=>nx7741, A1=>nx7401, B0=>nx7769);
   i8_ix75 : dffr port map ( Q=>i8_nx74, QB=>OPEN, D=>nx2, CLK=>CLK, R=>nx98
   );
   ix99 : nor02_2x port map ( Y=>nx98, A0=>nx3917, A1=>nx3919);
   ix3918 : nand02 port map ( Y=>nx3917, A0=>CNNIMGLOAD, A1=>nx7907);
   ix3920 : nand02 port map ( Y=>nx3919, A0=>nx7779, A1=>nx4083);
   i8_reg_start : dffs_ni port map ( Q=>OPEN, QB=>nx3921, D=>nx3293, CLK=>
      CLK, S=>nx588);
   ix3294 : nor02_2x port map ( Y=>nx3293, A0=>nx7775, A1=>nx3104);
   ix579 : nor02_2x port map ( Y=>nx3104, A0=>nx3925, A1=>nx7769);
   ix573 : nor02_2x port map ( Y=>nx572, A0=>nx3917, A1=>nx3928);
   ix3929 : nand02 port map ( Y=>nx3928, A0=>nx7775, A1=>nx3930);
   ix3284 : nor02_2x port map ( Y=>nx3283, A0=>nx3930, A1=>nx546);
   ix547 : nand03 port map ( Y=>nx546, A0=>nx3935, A1=>nx4181, A2=>nx3955);
   ix529 : nand03 port map ( Y=>nx528, A0=>nx7781, A1=>nx7911, A2=>
      i8_counterout2_3);
   ix3939 : nor02_2x port map ( Y=>nx3938, A0=>nx3940, A1=>nx4126);
   ix3208 : oai21 port map ( Y=>nx3207, A0=>nx3943, A1=>nx7785, B0=>nx4179);
   ix377 : nand02 port map ( Y=>nx376, A0=>nx3947, A1=>nx7737);
   ix3948 : nor02_2x port map ( Y=>nx3947, A0=>i8_reset2, A1=>nx7741);
   i8_ix97 : dffr port map ( Q=>i8_reset2, QB=>nx3925, D=>nx2, CLK=>CLK, R=>
      nx572);
   reg_i8_counterout2_0 : dff port map ( Q=>i8_counterout2_0, QB=>nx3940, D
      =>nx3207, CLK=>CLK);
   ix537 : nor02_2x port map ( Y=>nx536, A0=>nx3959, A1=>nx4093);
   ix3960 : nor02_2x port map ( Y=>nx3959, A0=>nx360, A1=>nx356);
   ix361 : nand04 port map ( Y=>nx360, A0=>nx3962, A1=>nx3979, A2=>nx4059, 
      A3=>i8_counterout1_0);
   ix3963 : nor02_2x port map ( Y=>nx3962, A0=>i8_counterout1_4, A1=>
      i8_counterout1_5);
   ix207 : oai22 port map ( Y=>nx206, A0=>nx3967, A1=>nx3969, B0=>nx3095, B1
      =>nx104);
   reg_i8_counterout1_4 : dff port map ( Q=>i8_counterout1_4, QB=>nx3967, D
      =>nx3157, CLK=>CLK);
   ix3970 : mux21 port map ( Y=>nx3969, A0=>nx7769, A1=>nx3093, S0=>nx7801);
   ix3972 : nor03_2x port map ( Y=>nx3971, A0=>nx7415, A1=>nx7741, A2=>
      nx7401);
   ix299 : nand04 port map ( Y=>nx298, A0=>nx3976, A1=>nx4083, A2=>
      loadingCNN, A3=>nx7775);
   ix3977 : oai21 port map ( Y=>nx3976, A0=>nx3093, A1=>nx282, B0=>nx3955);
   ix283 : nand03 port map ( Y=>nx282, A0=>nx3962, A1=>nx3979, A2=>nx4059);
   ix255 : oai22 port map ( Y=>nx254, A0=>nx3979, A1=>nx3985, B0=>nx3099, B1
      =>nx104);
   ix3986 : mux21 port map ( Y=>nx3985, A0=>nx7769, A1=>nx3097, S0=>nx7801);
   ix239 : nand04 port map ( Y=>nx3097, A0=>nx3988, A1=>nx4033, A2=>nx3967, 
      A3=>nx4050);
   ix3989 : nor03_2x port map ( Y=>nx3988, A0=>i8_counterout1_0, A1=>
      i8_counterout1_1, A2=>i8_counterout1_2);
   ix3198 : oai21 port map ( Y=>nx3197, A0=>nx3993, A1=>nx7803, B0=>nx4075);
   ix3994 : aoi322 port map ( Y=>nx3993, A0=>nx330, A1=>nx54, A2=>nx7413, B0
      =>nx3899, B1=>nx7799, C0=>i8_counterout1_1, C1=>nx340);
   ix331 : nand02 port map ( Y=>nx330, A0=>DataBus(14), A1=>DataBus(15));
   ix55 : inv01 port map ( Y=>nx54, A=>nx3541);
   ix341 : mux21 port map ( Y=>nx340, A0=>nx7413, A1=>nx3907, S0=>nx7799);
   ix4000 : nand02 port map ( Y=>nx3999, A0=>loadingCNN, A1=>nx316);
   ix317 : nand03 port map ( Y=>nx316, A0=>nx4002, A1=>i8_read2, A2=>nx7775
   );
   ix4003 : nand02 port map ( Y=>nx4002, A0=>nx7413, A1=>zed);
   ix541 : nor03_2x port map ( Y=>nx540, A0=>nx4007, A1=>nx3093, A2=>nx282);
   ix4008 : nand02 port map ( Y=>nx4007, A0=>i8_reset2, A1=>nx7413);
   i8_reg_read2 : dffs_ni port map ( Q=>i8_read2, QB=>nx3930, D=>nx3283, CLK
      =>CLK, S=>nx560);
   ix561 : nand03 port map ( Y=>nx560, A0=>nx546, A1=>nx4011, A2=>nx7775);
   ix4012 : nand04 port map ( Y=>nx4011, A0=>nx4013, A1=>nx4045, A2=>nx3541, 
      A3=>nx7395);
   ix167 : nand03 port map ( Y=>nx3092, A0=>nx3907, A1=>nx4016, A2=>nx4019);
   reg_i8_counterout1_1 : dff port map ( Q=>i8_counterout1_1, QB=>nx4016, D
      =>nx3197, CLK=>CLK);
   ix3138 : oai21 port map ( Y=>nx3137, A0=>nx4022, A1=>nx7803, B0=>nx4026);
   ix4023 : aoi322 port map ( Y=>nx4022, A0=>nx7413, A1=>DataBus(15), A2=>
      DataBus(14), B0=>nx3988, B1=>nx7799, C0=>i8_counterout1_2, C1=>nx152);
   reg_i8_counterout1_2 : dff port map ( Q=>i8_counterout1_2, QB=>nx4019, D
      =>nx3137, CLK=>CLK);
   ix153 : mux21 port map ( Y=>nx152, A0=>nx7413, A1=>nx3899, S0=>nx7799);
   ix4027 : oai21 port map ( Y=>nx4026, A0=>nx3917, A1=>nx4029, B0=>
      i8_counterout1_2);
   ix315 : oai21 port map ( Y=>nx314, A0=>nx7769, A1=>nx3955, B0=>i8_read2);
   ix183 : oai22 port map ( Y=>nx182, A0=>nx4033, A1=>nx4037, B0=>nx3093, B1
      =>nx104);
   ix4038 : mux21 port map ( Y=>nx4037, A0=>nx7769, A1=>nx3092, S0=>nx7799);
   ix105 : nand02 port map ( Y=>nx104, A0=>nx4041, A1=>nx7737);
   ix4042 : nor02_2x port map ( Y=>nx4041, A0=>nx7413, A1=>nx7741);
   reg_i8_counterout1_3 : dff port map ( Q=>i8_counterout1_3, QB=>nx4033, D
      =>nx3147, CLK=>CLK);
   ix4046 : nor03_2x port map ( Y=>nx4045, A0=>i8_counterout1_4, A1=>
      i8_counterout1_5, A2=>nx278);
   ix231 : oai22 port map ( Y=>nx230, A0=>nx4050, A1=>nx4053, B0=>nx3097, B1
      =>nx104);
   reg_i8_counterout1_5 : dff port map ( Q=>i8_counterout1_5, QB=>nx4050, D
      =>nx3167, CLK=>CLK);
   ix4054 : mux21 port map ( Y=>nx4053, A0=>nx7769, A1=>nx3095, S0=>nx7799);
   ix215 : nand04 port map ( Y=>nx3095, A0=>nx3899, A1=>nx4019, A2=>nx4033, 
      A3=>nx3967);
   ix279 : nand02 port map ( Y=>nx278, A0=>nx3979, A1=>nx4059);
   ix3188 : oai21 port map ( Y=>nx3187, A0=>nx4063, A1=>nx7803, B0=>nx4073);
   ix4064 : nor02_2x port map ( Y=>nx4063, A0=>nx268, A1=>nx110);
   ix269 : nor02_2x port map ( Y=>nx268, A0=>nx4066, A1=>nx104);
   reg_i8_counterout1_7 : dff port map ( Q=>i8_counterout1_7, QB=>nx4059, D
      =>nx3187, CLK=>CLK);
   ix111 : nor03_2x port map ( Y=>nx110, A0=>nx4059, A1=>nx7415, A2=>nx7799
   );
   ix4074 : oai21 port map ( Y=>nx4073, A0=>nx3917, A1=>nx4029, B0=>
      i8_counterout1_7);
   ix4076 : oai21 port map ( Y=>nx4075, A0=>nx3917, A1=>nx4029, B0=>
      i8_counterout1_1);
   ix263 : nand02 port map ( Y=>nx3099, A0=>nx4079, A1=>nx3979);
   i8_counterout1_6 : dff port map ( Q=>OPEN, QB=>nx3979, D=>nx3177, CLK=>
      CLK);
   i8_ix263 : dffsr_ni port map ( Q=>EnableReadingFromCPU2, QB=>nx4083, D=>
      DecompressedData1(255), CLK=>CLK, S=>nx610, R=>nx622);
   ix623 : nor02ii port map ( Y=>nx622, A0=>nx610, A1=>nx618);
   ix619 : oai221 port map ( Y=>nx618, A0=>zed, A1=>nx362, B0=>DataBus(14), 
      B1=>DataBus(15), C0=>nx7775);
   ix363 : nand04 port map ( Y=>nx362, A0=>nx4045, A1=>i8_counterout1_0, A2
      =>nx4090, A3=>nx4016);
   ix4091 : nor02_2x port map ( Y=>nx4090, A0=>i8_counterout1_2, A1=>
      i8_counterout1_3);
   ix357 : nand03 port map ( Y=>nx356, A0=>nx4019, A1=>nx4033, A2=>nx4016);
   ix4094 : nor02_2x port map ( Y=>nx4093, A0=>nx532, A1=>nx514);
   ix533 : nand04 port map ( Y=>nx532, A0=>nx7781, A1=>nx7911, A2=>
      i8_counterout2_3, A3=>i8_counterout2_4);
   ix3228 : inv01 port map ( Y=>nx3227, A=>nx4100);
   ix4101 : nor02_2x port map ( Y=>nx4100, A0=>nx3223, A1=>nx3225);
   ix3224 : nor02_2x port map ( Y=>nx3223, A0=>nx7961, A1=>nx7419);
   reg_i8_counterout2_2 : dff port map ( Q=>i8_counterout2_2, QB=>OPEN, D=>
      nx3227, CLK=>CLK);
   ix371 : nand03 port map ( Y=>nx370, A0=>nx7811, A1=>nx7395, A2=>nx7777);
   ix4108 : nand02 port map ( Y=>nx4107, A0=>i8_reset2, A1=>zed);
   ix3226 : aoi32 port map ( Y=>nx3225, A0=>nx7811, A1=>nx7395, A2=>nx7777, 
      B0=>nx4111, B1=>nx3102);
   ix4112 : nor03_2x port map ( Y=>nx4111, A0=>nx408, A1=>nx7427, A2=>nx7401
   );
   ix409 : nor02_2x port map ( Y=>nx408, A0=>nx7961, A1=>nx7813);
   ix4115 : nor02_2x port map ( Y=>nx4114, A0=>i8_counterout2_0, A1=>
      i8_counterout2_1);
   reg_i8_counterout2_1 : dff port map ( Q=>i8_counterout2_1, QB=>nx4126, D
      =>nx3217, CLK=>CLK);
   ix3218 : oai21 port map ( Y=>nx3217, A0=>nx4119, A1=>nx7785, B0=>nx4124);
   ix4120 : nor03_2x port map ( Y=>nx4119, A0=>nx396, A1=>nx7427, A2=>nx7401
   );
   ix375 : nand02 port map ( Y=>nx374, A0=>nx3925, A1=>CNNIMGLOAD);
   ix4125 : nand04 port map ( Y=>nx4124, A0=>i8_counterout2_1, A1=>nx7811, 
      A2=>nx7395, A3=>nx7777);
   ix423 : nand03 port map ( Y=>nx3102, A0=>nx3940, A1=>nx4126, A2=>nx7961);
   ix3238 : inv01 port map ( Y=>nx3237, A=>nx4131);
   ix4132 : nor02_2x port map ( Y=>nx4131, A0=>nx3233, A1=>nx3235);
   ix3234 : nor02_2x port map ( Y=>nx3233, A0=>nx7815, A1=>nx7419);
   reg_i8_counterout2_3 : dff port map ( Q=>i8_counterout2_3, QB=>OPEN, D=>
      nx3237, CLK=>CLK);
   ix3236 : aoi32 port map ( Y=>nx3235, A0=>nx7811, A1=>nx7395, A2=>nx7777, 
      B0=>nx4138, B1=>nx3101);
   ix4139 : nor03_2x port map ( Y=>nx4138, A0=>nx424, A1=>nx7427, A2=>nx7401
   );
   ix425 : nor02_2x port map ( Y=>nx424, A0=>nx7815, A1=>nx4141);
   ix4142 : nor03_2x port map ( Y=>nx4141, A0=>i8_counterout2_0, A1=>
      i8_counterout2_1, A2=>nx7911);
   ix439 : nand03 port map ( Y=>nx3101, A0=>nx7813, A1=>nx7961, A2=>nx7815);
   reg_i8_counterout2_4 : dff port map ( Q=>i8_counterout2_4, QB=>nx4151, D
      =>nx3247, CLK=>CLK);
   ix3248 : inv01 port map ( Y=>nx3247, A=>nx4148);
   ix4149 : aoi44 port map ( Y=>nx4148, A0=>i8_counterout2_4, A1=>nx7811, A2
      =>nx7395, A3=>nx7777, B0=>nx3947, B1=>nx7737, B2=>nx444, B3=>nx7419);
   ix515 : nand03 port map ( Y=>nx514, A0=>i8_counterout2_6, A1=>
      i8_counterout2_7, A2=>i8_counterout2_5);
   reg_i8_counterout2_6 : dff port map ( Q=>i8_counterout2_6, QB=>nx4167, D
      =>nx3267, CLK=>CLK);
   ix3268 : inv01 port map ( Y=>nx3267, A=>nx4155);
   ix4156 : aoi44 port map ( Y=>nx4155, A0=>i8_counterout2_6, A1=>nx7811, A2
      =>nx7395, A3=>nx7777, B0=>nx3947, B1=>nx7737, B2=>nx480, B3=>nx7419);
   ix459 : nand04 port map ( Y=>nx458, A0=>nx4141, A1=>nx7815, A2=>nx4151, 
      A3=>nx4159);
   ix3258 : inv01 port map ( Y=>nx3257, A=>nx4162);
   ix4163 : aoi44 port map ( Y=>nx4162, A0=>i8_counterout2_5, A1=>nx4107, A2
      =>nx7397, A3=>nx7777, B0=>nx3947, B1=>nx7737, B2=>nx464, B3=>nx7419);
   reg_i8_counterout2_5 : dff port map ( Q=>i8_counterout2_5, QB=>nx4159, D
      =>nx3257, CLK=>CLK);
   ix457 : nand04 port map ( Y=>nx3100, A0=>nx7813, A1=>nx7961, A2=>nx7815, 
      A3=>nx4151);
   reg_i8_counterout2_7 : dff port map ( Q=>i8_counterout2_7, QB=>nx4177, D
      =>nx3277, CLK=>CLK);
   ix3278 : inv01 port map ( Y=>nx3277, A=>nx4171);
   ix4172 : aoi44 port map ( Y=>nx4171, A0=>i8_counterout2_7, A1=>nx4107, A2
      =>nx7397, A3=>nx7779, B0=>nx494, B1=>nx3947, B2=>nx7739, B3=>nx7419);
   ix4180 : nand04 port map ( Y=>nx4179, A0=>i8_counterout2_0, A1=>nx7811, 
      A2=>nx7397, A3=>nx7779);
   ix4182 : nor03_2x port map ( Y=>nx4181, A0=>nx4167, A1=>nx4177, A2=>
      nx4159);
   ix589 : nor02_2x port map ( Y=>nx588, A0=>i8_loadenableD, A1=>nx3917);
   i8_reg_loadenableD : dff port map ( Q=>i8_loadenableD, QB=>OPEN, D=>
      loadingCNN, CLK=>CLK);
   ix4189 : nand02 port map ( Y=>nx4188, A0=>nx4191, A1=>nx7415);
   ix4192 : inv01 port map ( Y=>nx4191, A=>DataBus(14));
   ix129 : nor03_2x port map ( Y=>nx128, A0=>i8_counterout1_0, A1=>nx102, A2
      =>nx7401);
   ix103 : nand02 port map ( Y=>nx102, A0=>nx7771, A1=>CNNIMGLOAD);
   ix4197 : oai21 port map ( Y=>nx4196, A0=>nx3917, A1=>nx4029, B0=>
      i8_counterout1_0);
   ix603 : oai21 port map ( Y=>nx602, A0=>zed, A1=>nx362, B0=>nx54);
   ix3484 : nor02_2x port map ( Y=>nx3483, A0=>nx4203, A1=>nx1154);
   i7_reg_read1 : dffs_ni port map ( Q=>EnableReadingFromCPU1, QB=>nx4203, D
      =>nx3483, CLK=>CLK, S=>nx1158);
   ix1159 : nand02 port map ( Y=>nx1158, A0=>nx1154, A1=>nx7823);
   ix1155 : nand04 port map ( Y=>nx1154, A0=>nx4207, A1=>nx4370, A2=>nx4447, 
      A3=>nx4277);
   ix4208 : nor03_2x port map ( Y=>nx4207, A0=>nx4209, A1=>i7_counterout1_1, 
      A2=>nx1130);
   ix3408 : oai21 port map ( Y=>nx3407, A0=>nx4212, A1=>nx7835, B0=>nx4517);
   ix4213 : nor02_2x port map ( Y=>nx4212, A0=>nx960, A1=>nx952);
   ix961 : oai21 port map ( Y=>nx960, A0=>nx4209, A1=>nx4215, B0=>nx4509);
   ix4216 : oai21 port map ( Y=>nx4215, A0=>CNNIMGLOAD, A1=>nx7401, B0=>
      nx4217);
   ix639 : nor03_2x port map ( Y=>nx638, A0=>CNNIMGLOAD, A1=>nx7957, A2=>
      nx4220);
   ix4221 : nand02 port map ( Y=>nx4220, A0=>nx7823, A1=>nx4203);
   ix3394 : nor02_2x port map ( Y=>nx3393, A0=>nx7819, A1=>nx836);
   ix837 : nor02_2x port map ( Y=>nx836, A0=>nx4217, A1=>nx4227);
   ix831 : nor03_2x port map ( Y=>nx830, A0=>CNNIMGLOAD, A1=>nx7957, A2=>
      nx4231);
   ix4232 : nand02 port map ( Y=>nx4231, A0=>nx7819, A1=>nx4233);
   ix3384 : nor02_2x port map ( Y=>nx3383, A0=>nx4233, A1=>nx814);
   ix815 : nand04 port map ( Y=>nx814, A0=>nx4237, A1=>nx4281, A2=>nx4343, 
      A3=>nx4277);
   ix4238 : nor03_2x port map ( Y=>nx4237, A0=>nx4239, A1=>nx4318, A2=>nx802
   );
   ix3328 : inv01 port map ( Y=>nx3327, A=>nx4243);
   ix4244 : aoi44 port map ( Y=>nx4243, A0=>i7_counterout2_2, A1=>nx7827, A2
      =>nx7392, A3=>nx7821, B0=>nx4301, B1=>nx7739, B2=>nx690, B3=>nx650);
   reg_i7_counterout2_2 : dff port map ( Q=>i7_counterout2_2, QB=>nx4239, D
      =>nx3327, CLK=>CLK);
   ix4247 : nand02 port map ( Y=>nx4246, A0=>i7_reset2, A1=>i7_tmp);
   i7_ix81 : dffr port map ( Q=>i7_reset2, QB=>nx4227, D=>nx2, CLK=>CLK, R=>
      nx830);
   ix1141 : nor02_2x port map ( Y=>nx1140, A0=>nx4251, A1=>nx4501);
   ix4252 : nor03_2x port map ( Y=>nx4251, A0=>nx1134, A1=>nx1130, A2=>
      nx1128);
   ix1135 : nand02 port map ( Y=>nx1134, A0=>i7_counterout1_0, A1=>nx4255);
   reg_i7_counterout1_0 : dff port map ( Q=>i7_counterout1_0, QB=>nx4209, D
      =>nx3407, CLK=>CLK);
   ix3418 : oai21 port map ( Y=>nx3417, A0=>nx4258, A1=>nx7833, B0=>nx4496);
   ix4259 : aoi322 port map ( Y=>nx4258, A0=>nx940, A1=>nx4263, A2=>nx7441, 
      B0=>nx4267, B1=>nx7829, C0=>i7_counterout1_1, C1=>nx974);
   ix941 : inv01 port map ( Y=>nx940, A=>nx4261);
   ix4262 : nor02_2x port map ( Y=>nx4261, A0=>DataBus(9), A1=>DataBus(8));
   ix4264 : nand02 port map ( Y=>nx4263, A0=>DataBus(8), A1=>DataBus(9));
   i7_ix59 : dffr port map ( Q=>OPEN, QB=>nx4217, D=>nx2, CLK=>CLK, R=>nx638
   );
   ix4268 : nor02_2x port map ( Y=>nx4267, A0=>i7_counterout1_0, A1=>
      i7_counterout1_1);
   reg_i7_counterout1_1 : dff port map ( Q=>i7_counterout1_1, QB=>nx4255, D
      =>nx3417, CLK=>CLK);
   ix4272 : nor03_2x port map ( Y=>nx4271, A0=>nx7441, A1=>CNNIMGLOAD, A2=>
      nx7403);
   ix975 : mux21 port map ( Y=>nx974, A0=>nx7441, A1=>nx4209, S0=>nx7829);
   ix4275 : oai21 port map ( Y=>nx4274, A0=>nx856, A1=>i7_start, B0=>
      loadingimg);
   ix857 : oai21 port map ( Y=>nx856, A0=>nx4217, A1=>nx4277, B0=>i7_read2);
   ix1149 : nor03_2x port map ( Y=>nx1148, A0=>nx812, A1=>nx4367, A2=>nx1138
   );
   ix813 : nand03 port map ( Y=>nx812, A0=>nx4237, A1=>nx4281, A2=>nx4343);
   ix4282 : nor02_2x port map ( Y=>nx4281, A0=>nx4283, A1=>nx4333);
   ix3348 : oai21 port map ( Y=>nx3347, A0=>nx4287, A1=>nx7839, B0=>nx4331);
   ix4288 : nor03_2x port map ( Y=>nx4287, A0=>nx724, A1=>nx7447, A2=>nx7403
   );
   reg_i7_counterout2_4 : dff port map ( Q=>i7_counterout2_4, QB=>nx4283, D
      =>nx3347, CLK=>CLK);
   ix719 : nand03 port map ( Y=>nx3111, A0=>nx7837, A1=>nx4239, A2=>nx4318);
   ix4294 : nor02_2x port map ( Y=>nx4293, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1);
   reg_i7_counterout2_0 : dff port map ( Q=>i7_counterout2_0, QB=>nx4309, D
      =>nx3307, CLK=>CLK);
   ix3308 : oai21 port map ( Y=>nx3307, A0=>nx4298, A1=>nx7839, B0=>nx4307);
   ix655 : nand02 port map ( Y=>nx654, A0=>nx4301, A1=>nx7739);
   ix4302 : nor02_2x port map ( Y=>nx4301, A0=>i7_reset2, A1=>CNNIMGLOAD);
   ix649 : oai21 port map ( Y=>nx648, A0=>nx4227, A1=>nx4277, B0=>nx7390);
   ix4308 : nand04 port map ( Y=>nx4307, A0=>i7_counterout2_0, A1=>nx7825, 
      A2=>nx7390, A3=>nx7819);
   reg_i7_counterout2_1 : dff port map ( Q=>i7_counterout2_1, QB=>nx4317, D
      =>nx3317, CLK=>CLK);
   ix3318 : oai21 port map ( Y=>nx3317, A0=>nx4312, A1=>nx7839, B0=>nx4315);
   ix4313 : nor04 port map ( Y=>nx4312, A0=>nx674, A1=>i7_reset2, A2=>
      CNNIMGLOAD, A3=>nx7403);
   ix4316 : nand04 port map ( Y=>nx4315, A0=>i7_counterout2_1, A1=>nx7825, 
      A2=>nx7390, A3=>nx7819);
   ix3338 : oai21 port map ( Y=>nx3337, A0=>nx4322, A1=>nx7839, B0=>nx4327);
   ix4323 : nor04 port map ( Y=>nx4322, A0=>nx708, A1=>i7_reset2, A2=>
      CNNIMGLOAD, A3=>nx7403);
   reg_i7_counterout2_3 : dff port map ( Q=>i7_counterout2_3, QB=>nx4318, D
      =>nx3337, CLK=>CLK);
   ix4328 : nand04 port map ( Y=>nx4327, A0=>i7_counterout2_3, A1=>nx7825, 
      A2=>nx7390, A3=>nx7819);
   ix4332 : nand04 port map ( Y=>nx4331, A0=>i7_counterout2_4, A1=>nx7825, 
      A2=>nx7390, A3=>nx7819);
   ix3358 : inv01 port map ( Y=>nx3357, A=>nx4336);
   ix4337 : aoi44 port map ( Y=>nx4336, A0=>i7_counterout2_5, A1=>nx7825, A2
      =>nx7390, A3=>nx7821, B0=>nx4301, B1=>nx7739, B2=>nx740, B3=>nx650);
   reg_i7_counterout2_5 : dff port map ( Q=>i7_counterout2_5, QB=>nx4333, D
      =>nx3357, CLK=>CLK);
   ix735 : nand04 port map ( Y=>nx3109, A0=>nx7837, A1=>nx4239, A2=>nx4318, 
      A3=>nx4283);
   ix651 : nand03 port map ( Y=>nx650, A0=>nx7825, A1=>nx7390, A2=>nx7821);
   ix4344 : nor02_2x port map ( Y=>nx4343, A0=>nx4345, A1=>nx4355);
   ix3368 : inv01 port map ( Y=>nx3367, A=>nx4348);
   ix4349 : aoi44 port map ( Y=>nx4348, A0=>i7_counterout2_6, A1=>nx7825, A2
      =>nx7392, A3=>nx7821, B0=>nx4301, B1=>nx7739, B2=>nx758, B3=>nx650);
   reg_i7_counterout2_6 : dff port map ( Q=>i7_counterout2_6, QB=>nx4345, D
      =>nx3367, CLK=>CLK);
   ix753 : nand04 port map ( Y=>nx3107, A0=>nx4353, A1=>nx4318, A2=>nx4283, 
      A3=>nx4333);
   ix4354 : nor03_2x port map ( Y=>nx4353, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1, A2=>i7_counterout2_2);
   ix3378 : inv01 port map ( Y=>nx3377, A=>nx4359);
   ix4360 : aoi44 port map ( Y=>nx4359, A0=>i7_counterout2_7, A1=>nx7827, A2
      =>nx7392, A3=>nx7821, B0=>nx4301, B1=>nx7739, B2=>nx772, B3=>nx650);
   reg_i7_counterout2_7 : dff port map ( Q=>i7_counterout2_7, QB=>nx4355, D
      =>nx3377, CLK=>CLK);
   ix4368 : nand02 port map ( Y=>nx4367, A0=>nx7441, A1=>i7_reset2);
   ix1139 : nand03 port map ( Y=>nx1138, A0=>nx4207, A1=>nx4370, A2=>nx4447
   );
   ix4371 : nor02_2x port map ( Y=>nx4370, A0=>i7_counterout1_4, A1=>
      i7_counterout1_5);
   ix3448 : oai21 port map ( Y=>nx3447, A0=>nx4374, A1=>nx7833, B0=>nx4430);
   ix4375 : aoi322 port map ( Y=>nx4374, A0=>nx894, A1=>nx4383, A2=>nx7441, 
      B0=>nx4386, B1=>nx7829, C0=>i7_counterout1_4, C1=>nx1034);
   ix895 : oai21 port map ( Y=>nx894, A0=>nx4377, A1=>nx4379, B0=>nx4381);
   ix4378 : inv02 port map ( Y=>nx4377, A=>DataBus(11));
   ix4380 : nand03 port map ( Y=>nx4379, A0=>DataBus(10), A1=>DataBus(8), A2
      =>DataBus(9));
   ix4382 : inv02 port map ( Y=>nx4381, A=>DataBus(12));
   ix1029 : nand03 port map ( Y=>nx3117, A0=>nx4267, A1=>nx4389, A2=>nx4409
   );
   ix3428 : oai21 port map ( Y=>nx3427, A0=>nx4393, A1=>nx7833, B0=>nx4403);
   ix4394 : aoi322 port map ( Y=>nx4393, A0=>nx926, A1=>nx4379, A2=>nx7441, 
      B0=>nx4399, B1=>nx7829, C0=>i7_counterout1_2, C1=>nx994);
   ix927 : nand02 port map ( Y=>nx926, A0=>nx4263, A1=>nx4397);
   ix4398 : inv01 port map ( Y=>nx4397, A=>DataBus(10));
   ix4400 : nor03_2x port map ( Y=>nx4399, A0=>i7_counterout1_0, A1=>
      i7_counterout1_1, A2=>i7_counterout1_2);
   reg_i7_counterout1_2 : dff port map ( Q=>i7_counterout1_2, QB=>nx4389, D
      =>nx3427, CLK=>CLK);
   ix995 : mux21 port map ( Y=>nx994, A0=>nx7441, A1=>nx4267, S0=>nx7829);
   ix4404 : oai21 port map ( Y=>nx4403, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_2);
   ix4406 : nand02 port map ( Y=>nx4405, A0=>nx7741, A1=>nx7907);
   ix3438 : oai21 port map ( Y=>nx3437, A0=>nx4413, A1=>nx7833, B0=>nx4425);
   ix4414 : aoi322 port map ( Y=>nx4413, A0=>nx912, A1=>nx4417, A2=>nx7443, 
      B0=>nx4419, B1=>nx7829, C0=>i7_counterout1_3, C1=>nx1014);
   ix913 : oai21 port map ( Y=>nx912, A0=>nx4397, A1=>nx4263, B0=>nx4377);
   ix4418 : nand04 port map ( Y=>nx4417, A0=>DataBus(11), A1=>DataBus(10), 
      A2=>DataBus(8), A3=>DataBus(9));
   ix1009 : nand03 port map ( Y=>nx3118, A0=>nx4209, A1=>nx4255, A2=>nx4389
   );
   reg_i7_counterout1_3 : dff port map ( Q=>i7_counterout1_3, QB=>nx4409, D
      =>nx3437, CLK=>CLK);
   ix1015 : mux21 port map ( Y=>nx1014, A0=>nx7443, A1=>nx4399, S0=>nx7829);
   ix4426 : oai21 port map ( Y=>nx4425, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_3);
   reg_i7_counterout1_4 : dff port map ( Q=>i7_counterout1_4, QB=>nx4427, D
      =>nx3447, CLK=>CLK);
   ix1035 : mux21 port map ( Y=>nx1034, A0=>nx7443, A1=>nx4419, S0=>nx7831);
   ix4431 : oai21 port map ( Y=>nx4430, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_4);
   ix3458 : oai21 port map ( Y=>nx3457, A0=>nx4434, A1=>nx7833, B0=>nx4445);
   ix4435 : aoi222 port map ( Y=>nx4434, A0=>nx1058, A1=>nx7443, B0=>nx4437, 
      B1=>nx7831, C0=>i7_counterout1_5, C1=>nx1054);
   ix1059 : xnor2 port map ( Y=>nx1058, A0=>DataBus(13), A1=>nx4383);
   ix1049 : nand04 port map ( Y=>nx3116, A0=>nx4267, A1=>nx4389, A2=>nx4409, 
      A3=>nx4427);
   reg_i7_counterout1_5 : dff port map ( Q=>i7_counterout1_5, QB=>nx4441, D
      =>nx3457, CLK=>CLK);
   ix1055 : mux21 port map ( Y=>nx1054, A0=>nx7443, A1=>nx4386, S0=>nx7831);
   ix4446 : oai21 port map ( Y=>nx4445, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_5);
   ix4448 : nor02_2x port map ( Y=>nx4447, A0=>i7_counterout1_6, A1=>
      i7_counterout1_7);
   ix3468 : oai21 port map ( Y=>nx3467, A0=>nx4453, A1=>nx7833, B0=>nx4469);
   ix4454 : aoi222 port map ( Y=>nx4453, A0=>nx1084, A1=>nx7443, B0=>nx4462, 
      B1=>nx7831, C0=>i7_counterout1_6, C1=>nx1078);
   ix1085 : inv01 port map ( Y=>nx1084, A=>nx4457);
   ix4458 : xnor2 port map ( Y=>nx4457, A0=>DataBus(14), A1=>nx1082);
   ix1083 : nor03_2x port map ( Y=>nx1082, A0=>nx4460, A1=>nx4381, A2=>
      nx4417);
   ix4461 : inv01 port map ( Y=>nx4460, A=>DataBus(13));
   ix1073 : nand04 port map ( Y=>nx3115, A0=>nx4399, A1=>nx4409, A2=>nx4427, 
      A3=>nx4441);
   reg_i7_counterout1_6 : dff port map ( Q=>i7_counterout1_6, QB=>nx4465, D
      =>nx3467, CLK=>CLK);
   ix1079 : mux21 port map ( Y=>nx1078, A0=>nx7443, A1=>nx4437, S0=>nx7831);
   ix4470 : oai21 port map ( Y=>nx4469, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_6);
   reg_i7_counterout1_7 : dff port map ( Q=>i7_counterout1_7, QB=>nx4487, D
      =>nx3477, CLK=>CLK);
   ix3478 : oai21 port map ( Y=>nx3477, A0=>nx4475, A1=>nx7833, B0=>nx4485);
   ix4476 : aoi222 port map ( Y=>nx4475, A0=>nx1110, A1=>nx7445, B0=>nx1100, 
      B1=>nx7831, C0=>i7_counterout1_7, C1=>nx874);
   ix1111 : xnor2 port map ( Y=>nx1110, A0=>DataBus(15), A1=>nx4479);
   ix4480 : nand02 port map ( Y=>nx4479, A0=>DataBus(14), A1=>nx1082);
   ix875 : nor02_2x port map ( Y=>nx874, A0=>nx7445, A1=>nx7831);
   ix4486 : oai21 port map ( Y=>nx4485, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_7);
   i7_reg_read2 : dffs_ni port map ( Q=>i7_read2, QB=>nx4233, D=>nx3383, CLK
      =>CLK, S=>nx818);
   ix819 : nand02 port map ( Y=>nx818, A0=>nx814, A1=>nx7821);
   i7_reg_start : dffs_ni port map ( Q=>i7_start, QB=>OPEN, D=>nx3393, CLK=>
      CLK, S=>nx846);
   ix847 : nor03_2x port map ( Y=>nx846, A0=>i7_loadenableD, A1=>CNNIMGLOAD, 
      A2=>nx7957);
   i7_reg_loadenableD : dff port map ( Q=>i7_loadenableD, QB=>OPEN, D=>
      loadingimg, CLK=>CLK);
   ix4497 : oai21 port map ( Y=>nx4496, A0=>nx7843, A1=>nx7847, B0=>
      i7_counterout1_1);
   ix1131 : nand02 port map ( Y=>nx1130, A0=>nx4389, A1=>nx4409);
   ix1129 : nand03 port map ( Y=>nx1128, A0=>nx4370, A1=>nx4465, A2=>nx4487
   );
   ix4502 : nor03_2x port map ( Y=>nx4501, A0=>nx808, A1=>nx802, A2=>nx796);
   ix809 : nand02 port map ( Y=>nx808, A0=>i7_counterout2_2, A1=>
      i7_counterout2_3);
   ix803 : nand02 port map ( Y=>nx802, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1);
   ix797 : nand03 port map ( Y=>nx796, A0=>nx4281, A1=>i7_counterout2_6, A2
      =>i7_counterout2_7);
   ix4510 : nand02 port map ( Y=>nx4509, A0=>nx4511, A1=>nx7445);
   ix4512 : inv01 port map ( Y=>nx4511, A=>DataBus(8));
   ix953 : nor03_2x port map ( Y=>nx952, A0=>i7_counterout1_0, A1=>nx862, A2
      =>nx7403);
   ix863 : nand02 port map ( Y=>nx862, A0=>nx4217, A1=>nx7741);
   ix4518 : oai21 port map ( Y=>nx4517, A0=>nx7845, A1=>nx7849, B0=>
      i7_counterout1_0);
   ix2123 : nor02ii port map ( Y=>nx2122, A0=>nx7537, A1=>nx7455);
   ix2109 : nand02 port map ( Y=>nx2108, A0=>nx4522, A1=>nx7853);
   ix4523 : nand04 port map ( Y=>nx4522, A0=>nx4525, A1=>nx7765, A2=>nx7435, 
      A3=>nx7813);
   ix4526 : nor02_2x port map ( Y=>nx4525, A0=>nx7911, A1=>i8_counterout2_3
   );
   ix1189 : nor02_2x port map ( Y=>nx1188, A0=>nx4532, A1=>nx7785);
   ix4533 : inv01 port map ( Y=>nx4532, A=>DataBus(0));
   ix2119 : nand02 port map ( Y=>nx2118, A0=>nx4535, A1=>nx4537);
   ix4536 : nand03 port map ( Y=>nx4535, A0=>nx7813, A1=>nx7419, A2=>nx4525
   );
   ix4538 : nor03_2x port map ( Y=>nx4537, A0=>nx2106, A1=>nx7427, A2=>
      nx7403);
   ix2107 : nor02_2x port map ( Y=>nx2106, A0=>nx2098, A1=>nx4542);
   ix2099 : nand02 port map ( Y=>nx2098, A0=>nx7961, A1=>nx7815);
   ix4543 : nand03 port map ( Y=>nx4542, A0=>nx7765, A1=>nx7435, A2=>nx7813
   );
   ix2149 : nor02ii port map ( Y=>nx2148, A0=>nx7537, A1=>nx7459);
   ix1203 : nor02_2x port map ( Y=>nx1202, A0=>nx4547, A1=>nx7785);
   ix4548 : inv01 port map ( Y=>nx4547, A=>DataBus(1));
   ix2175 : nor02ii port map ( Y=>nx2174, A0=>nx7537, A1=>nx7463);
   ix1217 : nor02_2x port map ( Y=>nx1216, A0=>nx4553, A1=>nx7785);
   ix4554 : inv01 port map ( Y=>nx4553, A=>DataBus(2));
   ix2201 : nor02ii port map ( Y=>nx2200, A0=>nx7537, A1=>nx7467);
   ix1231 : nor02_2x port map ( Y=>nx1230, A0=>nx4558, A1=>nx7785);
   ix4559 : inv01 port map ( Y=>nx4558, A=>DataBus(3));
   ix2227 : nor02ii port map ( Y=>nx2226, A0=>nx7537, A1=>nx7471);
   ix1245 : nor02_2x port map ( Y=>nx1244, A0=>nx4565, A1=>nx7785);
   ix4566 : inv01 port map ( Y=>nx4565, A=>DataBus(4));
   ix2253 : nor02ii port map ( Y=>nx2252, A0=>nx7537, A1=>nx7475);
   ix1259 : nor02_2x port map ( Y=>nx1258, A0=>nx4570, A1=>nx7787);
   ix4571 : inv01 port map ( Y=>nx4570, A=>DataBus(5));
   ix2279 : nor02ii port map ( Y=>nx2278, A0=>nx7537, A1=>nx7479);
   ix1273 : nor02_2x port map ( Y=>nx1272, A0=>nx4577, A1=>nx7787);
   ix4578 : inv01 port map ( Y=>nx4577, A=>DataBus(6));
   ix2305 : nor02ii port map ( Y=>nx2304, A0=>nx2108, A1=>nx7483);
   ix1287 : nor02_2x port map ( Y=>nx1286, A0=>nx4582, A1=>nx7787);
   ix4583 : inv01 port map ( Y=>nx4582, A=>DataBus(7));
   ix2335 : nor02ii port map ( Y=>nx2334, A0=>nx2108, A1=>nx7487);
   ix1301 : nor02_2x port map ( Y=>nx1300, A0=>nx4511, A1=>nx7787);
   ix2359 : nor02ii port map ( Y=>nx2358, A0=>nx2108, A1=>nx7491);
   ix1315 : nor02_2x port map ( Y=>nx1314, A0=>nx4592, A1=>nx7787);
   ix4593 : inv01 port map ( Y=>nx4592, A=>DataBus(9));
   ix2383 : nor02ii port map ( Y=>nx2382, A0=>nx2108, A1=>nx7495);
   ix1329 : nor02_2x port map ( Y=>nx1328, A0=>nx4397, A1=>nx7787);
   ix2407 : nor02ii port map ( Y=>nx2406, A0=>nx2108, A1=>nx7499);
   ix1343 : nor02_2x port map ( Y=>nx1342, A0=>nx4377, A1=>nx7787);
   ix2431 : nor02ii port map ( Y=>nx2430, A0=>nx2108, A1=>nx7503);
   ix1357 : nor02_2x port map ( Y=>nx1356, A0=>nx4381, A1=>nx7789);
   i8_r1_lat_q_13 : latch port map ( Q=>DecompressedData2(15), D=>nx2444, 
      CLK=>nx7541);
   ix2445 : nor02ii port map ( Y=>nx2444, A0=>nx2108, A1=>nx7507);
   ix1371 : nor02_2x port map ( Y=>nx1370, A0=>nx4460, A1=>nx7789);
   ix2525 : nor02ii port map ( Y=>nx2524, A0=>nx7575, A1=>nx7455);
   ix2515 : nand02 port map ( Y=>nx2514, A0=>nx4613, A1=>nx7853);
   ix4614 : nand04 port map ( Y=>nx4613, A0=>nx4525, A1=>nx7765, A2=>nx7435, 
      A3=>nx7863);
   ix4616 : nor02_2x port map ( Y=>nx4615, A0=>nx3940, A1=>i8_counterout2_1
   );
   ix2521 : nand02 port map ( Y=>nx2520, A0=>nx4618, A1=>nx4621);
   ix4619 : nand03 port map ( Y=>nx4618, A0=>nx7863, A1=>nx7421, A2=>nx4525
   );
   ix4622 : nor03_2x port map ( Y=>nx4621, A0=>nx2512, A1=>nx7427, A2=>
      nx7405);
   ix2513 : nor02_2x port map ( Y=>nx2512, A0=>nx2098, A1=>nx4625);
   ix4626 : nand03 port map ( Y=>nx4625, A0=>nx7765, A1=>nx7435, A2=>nx7863
   );
   ix2549 : nor02ii port map ( Y=>nx2548, A0=>nx7575, A1=>nx7459);
   ix2573 : nor02ii port map ( Y=>nx2572, A0=>nx7575, A1=>nx7463);
   ix2597 : nor02ii port map ( Y=>nx2596, A0=>nx7575, A1=>nx7467);
   ix2621 : nor02ii port map ( Y=>nx2620, A0=>nx7575, A1=>nx7471);
   ix2645 : nor02ii port map ( Y=>nx2644, A0=>nx7575, A1=>nx7475);
   ix2669 : nor02ii port map ( Y=>nx2668, A0=>nx7575, A1=>nx7479);
   ix2693 : nor02ii port map ( Y=>nx2692, A0=>nx2514, A1=>nx7483);
   ix2723 : nor02ii port map ( Y=>nx2722, A0=>nx2514, A1=>nx7487);
   ix2747 : nor02ii port map ( Y=>nx2746, A0=>nx2514, A1=>nx7491);
   ix2771 : nor02ii port map ( Y=>nx2770, A0=>nx2514, A1=>nx7495);
   ix2795 : nor02ii port map ( Y=>nx2794, A0=>nx2514, A1=>nx7499);
   ix2819 : nor02ii port map ( Y=>nx2818, A0=>nx2514, A1=>nx7503);
   i8_r2_lat_q_13 : latch port map ( Q=>DecompressedData2(31), D=>nx2832, 
      CLK=>nx7579);
   ix2833 : nor02ii port map ( Y=>nx2832, A0=>nx2514, A1=>nx7507);
   ix2915 : nor02ii port map ( Y=>nx2914, A0=>nx7587, A1=>nx7455);
   ix2905 : nand02 port map ( Y=>nx2904, A0=>nx4663, A1=>nx7853);
   ix4664 : nand04 port map ( Y=>nx4663, A0=>nx4525, A1=>nx7765, A2=>nx7435, 
      A3=>nx7865);
   ix4666 : nor02_2x port map ( Y=>nx4665, A0=>i8_counterout2_0, A1=>nx4126
   );
   ix2911 : nand02 port map ( Y=>nx2910, A0=>nx4668, A1=>nx4670);
   ix4669 : nand03 port map ( Y=>nx4668, A0=>nx7865, A1=>nx7421, A2=>nx4525
   );
   ix4671 : nor03_2x port map ( Y=>nx4670, A0=>nx2902, A1=>nx7427, A2=>
      nx7405);
   ix2903 : nor02_2x port map ( Y=>nx2902, A0=>nx2098, A1=>nx4673);
   ix4674 : nand03 port map ( Y=>nx4673, A0=>nx7765, A1=>nx7435, A2=>nx7865
   );
   ix2939 : nor02ii port map ( Y=>nx2938, A0=>nx7587, A1=>nx7459);
   ix2963 : nor02ii port map ( Y=>nx2962, A0=>nx7587, A1=>nx7463);
   ix2987 : nor02ii port map ( Y=>nx2986, A0=>nx7587, A1=>nx7467);
   ix3011 : nor02ii port map ( Y=>nx3010, A0=>nx7587, A1=>nx7471);
   ix3035 : nor02ii port map ( Y=>nx3034, A0=>nx7587, A1=>nx7475);
   ix3059 : nor02ii port map ( Y=>nx3058, A0=>nx7587, A1=>nx7479);
   ix3083 : nor02ii port map ( Y=>nx3082, A0=>nx2904, A1=>nx7483);
   ix3113 : nor02ii port map ( Y=>nx3112, A0=>nx2904, A1=>nx7487);
   ix3137 : nor02ii port map ( Y=>nx3136, A0=>nx2904, A1=>nx7491);
   ix3161 : nor02ii port map ( Y=>nx3160, A0=>nx2904, A1=>nx7495);
   ix3185 : nor02ii port map ( Y=>nx3184, A0=>nx2904, A1=>nx7499);
   ix3209 : nor02ii port map ( Y=>nx3208, A0=>nx2904, A1=>nx7503);
   i8_r3_lat_q_13 : latch port map ( Q=>DecompressedData2(47), D=>nx3222, 
      CLK=>nx7591);
   ix3223 : nor02ii port map ( Y=>nx3222, A0=>nx2904, A1=>nx7507);
   ix3303 : nor02ii port map ( Y=>nx3302, A0=>nx7599, A1=>nx7455);
   ix3293 : nand02 port map ( Y=>nx3292, A0=>nx4711, A1=>nx7853);
   ix4712 : nand04 port map ( Y=>nx4711, A0=>nx4525, A1=>nx7767, A2=>nx7435, 
      A3=>nx7781);
   ix3299 : nand02 port map ( Y=>nx3298, A0=>nx4715, A1=>nx4717);
   ix4716 : nand03 port map ( Y=>nx4715, A0=>nx7781, A1=>nx7421, A2=>nx4525
   );
   ix4718 : nor03_2x port map ( Y=>nx4717, A0=>nx3290, A1=>nx7427, A2=>
      nx7405);
   ix3291 : nor02_2x port map ( Y=>nx3290, A0=>nx2098, A1=>nx4720);
   ix4721 : nand03 port map ( Y=>nx4720, A0=>nx7767, A1=>nx7437, A2=>nx7781
   );
   ix3327 : nor02ii port map ( Y=>nx3326, A0=>nx7599, A1=>nx7459);
   ix3351 : nor02ii port map ( Y=>nx3350, A0=>nx7599, A1=>nx7463);
   ix3375 : nor02ii port map ( Y=>nx3374, A0=>nx7599, A1=>nx7467);
   ix3399 : nor02ii port map ( Y=>nx3398, A0=>nx7599, A1=>nx7471);
   ix3423 : nor02ii port map ( Y=>nx3422, A0=>nx7599, A1=>nx7475);
   ix3447 : nor02ii port map ( Y=>nx3446, A0=>nx7599, A1=>nx7479);
   ix3471 : nor02ii port map ( Y=>nx3470, A0=>nx3292, A1=>nx7483);
   ix3501 : nor02ii port map ( Y=>nx3500, A0=>nx3292, A1=>nx7487);
   ix3525 : nor02ii port map ( Y=>nx3524, A0=>nx3292, A1=>nx7491);
   ix3549 : nor02ii port map ( Y=>nx3548, A0=>nx3292, A1=>nx7495);
   ix3573 : nor02ii port map ( Y=>nx3572, A0=>nx3292, A1=>nx7499);
   ix3597 : nor02ii port map ( Y=>nx3596, A0=>nx3292, A1=>nx7503);
   i8_r4_lat_q_13 : latch port map ( Q=>DecompressedData2(63), D=>nx3610, 
      CLK=>nx7603);
   ix3611 : nor02ii port map ( Y=>nx3610, A0=>nx3292, A1=>nx7507);
   ix3703 : nor02ii port map ( Y=>nx3702, A0=>nx7611, A1=>nx7455);
   ix3689 : nand02 port map ( Y=>nx3688, A0=>nx4757, A1=>nx7853);
   ix4758 : nand04 port map ( Y=>nx4757, A0=>nx4759, A1=>nx7767, A2=>nx7437, 
      A3=>nx7813);
   ix4760 : nor02_2x port map ( Y=>nx4759, A0=>nx7961, A1=>i8_counterout2_3
   );
   ix3699 : nand02 port map ( Y=>nx3698, A0=>nx4763, A1=>nx4765);
   ix4764 : nand03 port map ( Y=>nx4763, A0=>nx4114, A1=>nx7421, A2=>nx4759
   );
   ix4766 : nor03_2x port map ( Y=>nx4765, A0=>nx3686, A1=>nx7429, A2=>
      nx7405);
   ix3687 : nor02_2x port map ( Y=>nx3686, A0=>nx3682, A1=>nx4542);
   ix3683 : nand02 port map ( Y=>nx3682, A0=>nx7911, A1=>nx7815);
   ix3727 : nor02ii port map ( Y=>nx3726, A0=>nx7611, A1=>nx7459);
   ix3751 : nor02ii port map ( Y=>nx3750, A0=>nx7611, A1=>nx7463);
   ix3775 : nor02ii port map ( Y=>nx3774, A0=>nx7611, A1=>nx7467);
   ix3799 : nor02ii port map ( Y=>nx3798, A0=>nx7611, A1=>nx7471);
   ix3823 : nor02ii port map ( Y=>nx3822, A0=>nx7611, A1=>nx7475);
   ix3847 : nor02ii port map ( Y=>nx3846, A0=>nx7611, A1=>nx7479);
   ix3871 : nor02ii port map ( Y=>nx3870, A0=>nx3688, A1=>nx7483);
   ix3901 : nor02ii port map ( Y=>nx3900, A0=>nx3688, A1=>nx7487);
   ix3925 : nor02ii port map ( Y=>nx3924, A0=>nx3688, A1=>nx7491);
   ix3949 : nor02ii port map ( Y=>nx3948, A0=>nx3688, A1=>nx7495);
   ix3973 : nor02ii port map ( Y=>nx3972, A0=>nx3688, A1=>nx7499);
   ix3997 : nor02ii port map ( Y=>nx3996, A0=>nx3688, A1=>nx7503);
   i8_r5_lat_q_13 : latch port map ( Q=>DecompressedData2(79), D=>nx4010, 
      CLK=>nx7615);
   ix4011 : nor02ii port map ( Y=>nx4010, A0=>nx3688, A1=>nx7507);
   ix4087 : nor02ii port map ( Y=>nx4086, A0=>nx7623, A1=>nx7455);
   ix4077 : nand02 port map ( Y=>nx4076, A0=>nx4804, A1=>nx7853);
   ix4805 : nand04 port map ( Y=>nx4804, A0=>nx4759, A1=>nx7767, A2=>nx7437, 
      A3=>nx7863);
   ix4083 : nand02 port map ( Y=>nx4082, A0=>nx4807, A1=>nx4809);
   ix4808 : nand03 port map ( Y=>nx4807, A0=>nx7863, A1=>nx7421, A2=>nx4759
   );
   ix4810 : nor03_2x port map ( Y=>nx4809, A0=>nx4074, A1=>nx7429, A2=>
      nx7405);
   ix4075 : nor02_2x port map ( Y=>nx4074, A0=>nx3682, A1=>nx4625);
   ix4111 : nor02ii port map ( Y=>nx4110, A0=>nx7623, A1=>nx7459);
   ix4135 : nor02ii port map ( Y=>nx4134, A0=>nx7623, A1=>nx7463);
   ix4159 : nor02ii port map ( Y=>nx4158, A0=>nx7623, A1=>nx7467);
   ix4183 : nor02ii port map ( Y=>nx4182, A0=>nx7623, A1=>nx7471);
   ix4207 : nor02ii port map ( Y=>nx4206, A0=>nx7623, A1=>nx7475);
   ix4231 : nor02ii port map ( Y=>nx4230, A0=>nx7623, A1=>nx7479);
   ix4255 : nor02ii port map ( Y=>nx4254, A0=>nx4076, A1=>nx7483);
   ix4285 : nor02ii port map ( Y=>nx4284, A0=>nx4076, A1=>nx7487);
   ix4309 : nor02ii port map ( Y=>nx4308, A0=>nx4076, A1=>nx7491);
   ix4333 : nor02ii port map ( Y=>nx4332, A0=>nx4076, A1=>nx7495);
   ix4357 : nor02ii port map ( Y=>nx4356, A0=>nx4076, A1=>nx7499);
   ix4381 : nor02ii port map ( Y=>nx4380, A0=>nx4076, A1=>nx7503);
   i8_r6_lat_q_13 : latch port map ( Q=>DecompressedData2(95), D=>nx4394, 
      CLK=>nx7627);
   ix4395 : nor02ii port map ( Y=>nx4394, A0=>nx4076, A1=>nx7507);
   ix4481 : nor02ii port map ( Y=>nx4480, A0=>nx7643, A1=>nx7455);
   ix4471 : nand02 port map ( Y=>nx4470, A0=>nx4847, A1=>nx7853);
   ix4848 : nand04 port map ( Y=>nx4847, A0=>nx4759, A1=>nx7767, A2=>nx7437, 
      A3=>nx7865);
   ix4477 : nand02 port map ( Y=>nx4476, A0=>nx4851, A1=>nx4853);
   ix4852 : nand03 port map ( Y=>nx4851, A0=>nx7865, A1=>nx7421, A2=>nx4759
   );
   ix4854 : nor03_2x port map ( Y=>nx4853, A0=>nx4468, A1=>nx7429, A2=>
      nx7405);
   ix4469 : nor02_2x port map ( Y=>nx4468, A0=>nx3682, A1=>nx4673);
   ix4505 : nor02ii port map ( Y=>nx4504, A0=>nx7643, A1=>nx7459);
   ix4529 : nor02ii port map ( Y=>nx4528, A0=>nx7643, A1=>nx7463);
   ix4553 : nor02ii port map ( Y=>nx4552, A0=>nx7643, A1=>nx7467);
   ix4577 : nor02ii port map ( Y=>nx4576, A0=>nx7643, A1=>nx7471);
   ix4601 : nor02ii port map ( Y=>nx4600, A0=>nx7643, A1=>nx7475);
   ix4625 : nor02ii port map ( Y=>nx4624, A0=>nx7643, A1=>nx7479);
   ix4649 : nor02ii port map ( Y=>nx4648, A0=>nx4470, A1=>nx7483);
   ix4679 : nor02ii port map ( Y=>nx4678, A0=>nx4470, A1=>nx7487);
   ix4703 : nor02ii port map ( Y=>nx4702, A0=>nx4470, A1=>nx7491);
   ix4727 : nor02ii port map ( Y=>nx4726, A0=>nx4470, A1=>nx7495);
   ix4751 : nor02ii port map ( Y=>nx4750, A0=>nx4470, A1=>nx7499);
   ix4775 : nor02ii port map ( Y=>nx4774, A0=>nx4470, A1=>nx7503);
   i8_r7_lat_q_13 : latch port map ( Q=>DecompressedData2(111), D=>nx4788, 
      CLK=>nx7647);
   ix4789 : nor02ii port map ( Y=>nx4788, A0=>nx4470, A1=>nx7507);
   ix4865 : nor02ii port map ( Y=>nx4864, A0=>nx7655, A1=>nx7457);
   ix4855 : nand02 port map ( Y=>nx4854, A0=>nx4894, A1=>nx7855);
   ix4895 : nand04 port map ( Y=>nx4894, A0=>nx4759, A1=>nx7767, A2=>nx7437, 
      A3=>nx7781);
   ix4861 : nand02 port map ( Y=>nx4860, A0=>nx4897, A1=>nx4899);
   ix4898 : nand03 port map ( Y=>nx4897, A0=>nx7781, A1=>nx7421, A2=>nx4759
   );
   ix4900 : nor03_2x port map ( Y=>nx4899, A0=>nx4852, A1=>nx7429, A2=>
      nx7405);
   ix4853 : nor02_2x port map ( Y=>nx4852, A0=>nx3682, A1=>nx4720);
   ix4889 : nor02ii port map ( Y=>nx4888, A0=>nx7655, A1=>nx7461);
   ix4913 : nor02ii port map ( Y=>nx4912, A0=>nx7655, A1=>nx7465);
   ix4937 : nor02ii port map ( Y=>nx4936, A0=>nx7655, A1=>nx7469);
   ix4961 : nor02ii port map ( Y=>nx4960, A0=>nx7655, A1=>nx7473);
   ix4985 : nor02ii port map ( Y=>nx4984, A0=>nx7655, A1=>nx7477);
   ix5009 : nor02ii port map ( Y=>nx5008, A0=>nx7655, A1=>nx7481);
   ix5033 : nor02ii port map ( Y=>nx5032, A0=>nx4854, A1=>nx7485);
   ix5063 : nor02ii port map ( Y=>nx5062, A0=>nx4854, A1=>nx7489);
   ix5087 : nor02ii port map ( Y=>nx5086, A0=>nx4854, A1=>nx7493);
   ix5111 : nor02ii port map ( Y=>nx5110, A0=>nx4854, A1=>nx7497);
   ix5135 : nor02ii port map ( Y=>nx5134, A0=>nx4854, A1=>nx7501);
   ix5159 : nor02ii port map ( Y=>nx5158, A0=>nx4854, A1=>nx7505);
   i8_r8_lat_q_13 : latch port map ( Q=>DecompressedData2(127), D=>nx5172, 
      CLK=>nx7659);
   ix5173 : nor02ii port map ( Y=>nx5172, A0=>nx4854, A1=>nx7509);
   ix5263 : nor02ii port map ( Y=>nx5262, A0=>nx7667, A1=>nx7457);
   ix5249 : nand02 port map ( Y=>nx5248, A0=>nx4937, A1=>nx7855);
   ix4938 : nand04 port map ( Y=>nx4937, A0=>nx4939, A1=>nx7767, A2=>nx7437, 
      A3=>nx4114);
   ix4940 : nor02_2x port map ( Y=>nx4939, A0=>nx7911, A1=>nx7817);
   ix5259 : nand02 port map ( Y=>nx5258, A0=>nx4942, A1=>nx4945);
   ix4943 : nand03 port map ( Y=>nx4942, A0=>nx4114, A1=>nx7423, A2=>nx4939
   );
   ix4946 : nor03_2x port map ( Y=>nx4945, A0=>nx5246, A1=>nx7429, A2=>
      nx7407);
   ix5247 : nor02_2x port map ( Y=>nx5246, A0=>nx5242, A1=>nx4542);
   ix5243 : nand02 port map ( Y=>nx5242, A0=>nx7809, A1=>i8_counterout2_3);
   ix5287 : nor02ii port map ( Y=>nx5286, A0=>nx7667, A1=>nx7461);
   ix5311 : nor02ii port map ( Y=>nx5310, A0=>nx7667, A1=>nx7465);
   ix5335 : nor02ii port map ( Y=>nx5334, A0=>nx7667, A1=>nx7469);
   ix5359 : nor02ii port map ( Y=>nx5358, A0=>nx7667, A1=>nx7473);
   ix5383 : nor02ii port map ( Y=>nx5382, A0=>nx7667, A1=>nx7477);
   ix5407 : nor02ii port map ( Y=>nx5406, A0=>nx7667, A1=>nx7481);
   ix5431 : nor02ii port map ( Y=>nx5430, A0=>nx5248, A1=>nx7485);
   ix5461 : nor02ii port map ( Y=>nx5460, A0=>nx5248, A1=>nx7489);
   ix5485 : nor02ii port map ( Y=>nx5484, A0=>nx5248, A1=>nx7493);
   ix5509 : nor02ii port map ( Y=>nx5508, A0=>nx5248, A1=>nx7497);
   ix5533 : nor02ii port map ( Y=>nx5532, A0=>nx5248, A1=>nx7501);
   ix5557 : nor02ii port map ( Y=>nx5556, A0=>nx5248, A1=>nx7505);
   i8_r9_lat_q_13 : latch port map ( Q=>DecompressedData2(143), D=>nx5570, 
      CLK=>nx7671);
   ix5571 : nor02ii port map ( Y=>nx5570, A0=>nx5248, A1=>nx7509);
   ix5647 : nor02ii port map ( Y=>nx5646, A0=>nx7679, A1=>nx7457);
   ix5637 : nand02 port map ( Y=>nx5636, A0=>nx4985, A1=>nx7855);
   ix4986 : nand04 port map ( Y=>nx4985, A0=>nx4939, A1=>nx3895, A2=>nx7437, 
      A3=>nx7863);
   ix5643 : nand02 port map ( Y=>nx5642, A0=>nx4988, A1=>nx4990);
   ix4989 : nand03 port map ( Y=>nx4988, A0=>nx7863, A1=>nx7423, A2=>nx4939
   );
   ix4991 : nor03_2x port map ( Y=>nx4990, A0=>nx5634, A1=>nx7429, A2=>
      nx7407);
   ix5635 : nor02_2x port map ( Y=>nx5634, A0=>nx5242, A1=>nx4625);
   ix5671 : nor02ii port map ( Y=>nx5670, A0=>nx7679, A1=>nx7461);
   ix5695 : nor02ii port map ( Y=>nx5694, A0=>nx7679, A1=>nx7465);
   ix5719 : nor02ii port map ( Y=>nx5718, A0=>nx7679, A1=>nx7469);
   ix5743 : nor02ii port map ( Y=>nx5742, A0=>nx7679, A1=>nx7473);
   ix5767 : nor02ii port map ( Y=>nx5766, A0=>nx7679, A1=>nx7477);
   ix5791 : nor02ii port map ( Y=>nx5790, A0=>nx7679, A1=>nx7481);
   ix5815 : nor02ii port map ( Y=>nx5814, A0=>nx5636, A1=>nx7485);
   ix5845 : nor02ii port map ( Y=>nx5844, A0=>nx5636, A1=>nx7489);
   ix5869 : nor02ii port map ( Y=>nx5868, A0=>nx5636, A1=>nx7493);
   ix5893 : nor02ii port map ( Y=>nx5892, A0=>nx5636, A1=>nx7497);
   ix5917 : nor02ii port map ( Y=>nx5916, A0=>nx5636, A1=>nx7501);
   ix5941 : nor02ii port map ( Y=>nx5940, A0=>nx5636, A1=>nx7505);
   i8_r10_lat_q_13 : latch port map ( Q=>DecompressedData2(159), D=>nx5954, 
      CLK=>nx7683);
   ix5955 : nor02ii port map ( Y=>nx5954, A0=>nx5636, A1=>nx7509);
   ix6037 : nor02ii port map ( Y=>nx6036, A0=>nx7691, A1=>nx7457);
   ix6027 : nand02 port map ( Y=>nx6026, A0=>nx5029, A1=>nx7855);
   ix5030 : nand04 port map ( Y=>nx5029, A0=>nx4939, A1=>nx3895, A2=>nx7439, 
      A3=>nx7865);
   ix6033 : nand02 port map ( Y=>nx6032, A0=>nx5033, A1=>nx5035);
   ix5034 : nand03 port map ( Y=>nx5033, A0=>nx7865, A1=>nx7423, A2=>nx4939
   );
   ix5036 : nor03_2x port map ( Y=>nx5035, A0=>nx6024, A1=>nx7429, A2=>
      nx7407);
   ix6025 : nor02_2x port map ( Y=>nx6024, A0=>nx5242, A1=>nx4673);
   ix6061 : nor02ii port map ( Y=>nx6060, A0=>nx7691, A1=>nx7461);
   ix6085 : nor02ii port map ( Y=>nx6084, A0=>nx7691, A1=>nx7465);
   ix6109 : nor02ii port map ( Y=>nx6108, A0=>nx7691, A1=>nx7469);
   ix6133 : nor02ii port map ( Y=>nx6132, A0=>nx7691, A1=>nx7473);
   ix6157 : nor02ii port map ( Y=>nx6156, A0=>nx7691, A1=>nx7477);
   ix6181 : nor02ii port map ( Y=>nx6180, A0=>nx7691, A1=>nx7481);
   ix6205 : nor02ii port map ( Y=>nx6204, A0=>nx6026, A1=>nx7485);
   ix6235 : nor02ii port map ( Y=>nx6234, A0=>nx6026, A1=>nx7489);
   ix6259 : nor02ii port map ( Y=>nx6258, A0=>nx6026, A1=>nx7493);
   ix6283 : nor02ii port map ( Y=>nx6282, A0=>nx6026, A1=>nx7497);
   ix6307 : nor02ii port map ( Y=>nx6306, A0=>nx6026, A1=>nx7501);
   ix6331 : nor02ii port map ( Y=>nx6330, A0=>nx6026, A1=>nx7505);
   i8_r11_lat_q_13 : latch port map ( Q=>DecompressedData2(175), D=>nx6344, 
      CLK=>nx7695);
   ix6345 : nor02ii port map ( Y=>nx6344, A0=>nx6026, A1=>nx7509);
   ix6421 : nor02ii port map ( Y=>nx6420, A0=>nx7703, A1=>nx7457);
   ix6411 : nand02 port map ( Y=>nx6410, A0=>nx5075, A1=>nx7855);
   ix5076 : nand04 port map ( Y=>nx5075, A0=>nx4939, A1=>nx3895, A2=>nx7439, 
      A3=>nx3938);
   ix6417 : nand02 port map ( Y=>nx6416, A0=>nx5078, A1=>nx5080);
   ix5079 : nand03 port map ( Y=>nx5078, A0=>nx3938, A1=>nx7423, A2=>nx4939
   );
   ix5081 : nor03_2x port map ( Y=>nx5080, A0=>nx6408, A1=>nx7431, A2=>
      nx7407);
   ix6409 : nor02_2x port map ( Y=>nx6408, A0=>nx5242, A1=>nx4720);
   ix6445 : nor02ii port map ( Y=>nx6444, A0=>nx7703, A1=>nx7461);
   ix6469 : nor02ii port map ( Y=>nx6468, A0=>nx7703, A1=>nx7465);
   ix6493 : nor02ii port map ( Y=>nx6492, A0=>nx7703, A1=>nx7469);
   ix6517 : nor02ii port map ( Y=>nx6516, A0=>nx7703, A1=>nx7473);
   ix6541 : nor02ii port map ( Y=>nx6540, A0=>nx7703, A1=>nx7477);
   ix6565 : nor02ii port map ( Y=>nx6564, A0=>nx7703, A1=>nx7481);
   ix6589 : nor02ii port map ( Y=>nx6588, A0=>nx6410, A1=>nx7485);
   ix6619 : nor02ii port map ( Y=>nx6618, A0=>nx6410, A1=>nx7489);
   ix6643 : nor02ii port map ( Y=>nx6642, A0=>nx6410, A1=>nx7493);
   ix6667 : nor02ii port map ( Y=>nx6666, A0=>nx6410, A1=>nx7497);
   ix6691 : nor02ii port map ( Y=>nx6690, A0=>nx6410, A1=>nx7501);
   ix6715 : nor02ii port map ( Y=>nx6714, A0=>nx6410, A1=>nx7505);
   i8_r12_lat_q_13 : latch port map ( Q=>DecompressedData2(191), D=>nx6728, 
      CLK=>nx7707);
   ix6729 : nor02ii port map ( Y=>nx6728, A0=>nx6410, A1=>nx7509);
   ix6813 : nor02ii port map ( Y=>nx6812, A0=>nx7715, A1=>nx7457);
   ix6803 : nand02 port map ( Y=>nx6802, A0=>nx5119, A1=>nx7855);
   ix5120 : nand04 port map ( Y=>nx5119, A0=>nx5121, A1=>nx3895, A2=>nx7439, 
      A3=>nx4114);
   ix5122 : nor02_2x port map ( Y=>nx5121, A0=>nx7809, A1=>nx7817);
   ix6809 : nand02 port map ( Y=>nx6808, A0=>nx5124, A1=>nx5126);
   ix5125 : nand03 port map ( Y=>nx5124, A0=>nx4114, A1=>nx5121, A2=>nx7423
   );
   ix5127 : nor03_2x port map ( Y=>nx5126, A0=>nx6800, A1=>nx7431, A2=>
      nx7407);
   ix6801 : nor02_2x port map ( Y=>nx6800, A0=>nx520, A1=>nx4542);
   ix521 : nand02 port map ( Y=>nx520, A0=>nx7911, A1=>i8_counterout2_3);
   ix6837 : nor02ii port map ( Y=>nx6836, A0=>nx7715, A1=>nx7461);
   ix6861 : nor02ii port map ( Y=>nx6860, A0=>nx7715, A1=>nx7465);
   ix6885 : nor02ii port map ( Y=>nx6884, A0=>nx7715, A1=>nx7469);
   ix6909 : nor02ii port map ( Y=>nx6908, A0=>nx7715, A1=>nx7473);
   ix6933 : nor02ii port map ( Y=>nx6932, A0=>nx7715, A1=>nx7477);
   ix6957 : nor02ii port map ( Y=>nx6956, A0=>nx7715, A1=>nx7481);
   ix6981 : nor02ii port map ( Y=>nx6980, A0=>nx6802, A1=>nx7485);
   ix7011 : nor02ii port map ( Y=>nx7010, A0=>nx6802, A1=>nx7489);
   ix7035 : nor02ii port map ( Y=>nx7034, A0=>nx6802, A1=>nx7493);
   ix7059 : nor02ii port map ( Y=>nx7058, A0=>nx6802, A1=>nx7497);
   ix7083 : nor02ii port map ( Y=>nx7082, A0=>nx6802, A1=>nx7501);
   ix7107 : nor02ii port map ( Y=>nx7106, A0=>nx6802, A1=>nx7505);
   i8_r13_lat_q_13 : latch port map ( Q=>DecompressedData2(207), D=>nx7120, 
      CLK=>nx7719);
   ix7121 : nor02ii port map ( Y=>nx7120, A0=>nx6802, A1=>nx7509);
   ix7197 : nor02ii port map ( Y=>nx7196, A0=>nx7727, A1=>nx7457);
   ix7187 : nand02 port map ( Y=>nx7186, A0=>nx5165, A1=>nx7855);
   ix5166 : nand04 port map ( Y=>nx5165, A0=>nx5121, A1=>nx3895, A2=>nx7439, 
      A3=>nx4615);
   ix7193 : nand02 port map ( Y=>nx7192, A0=>nx5169, A1=>nx5171);
   ix5170 : nand03 port map ( Y=>nx5169, A0=>nx4615, A1=>nx5121, A2=>nx7423
   );
   ix5172 : nor03_2x port map ( Y=>nx5171, A0=>nx7184, A1=>nx7431, A2=>
      nx7407);
   ix7185 : nor02_2x port map ( Y=>nx7184, A0=>nx520, A1=>nx4625);
   ix7221 : nor02ii port map ( Y=>nx7220, A0=>nx7727, A1=>nx7461);
   ix7245 : nor02ii port map ( Y=>nx7244, A0=>nx7727, A1=>nx7465);
   ix7269 : nor02ii port map ( Y=>nx7268, A0=>nx7727, A1=>nx7469);
   ix7293 : nor02ii port map ( Y=>nx7292, A0=>nx7727, A1=>nx7473);
   ix7317 : nor02ii port map ( Y=>nx7316, A0=>nx7727, A1=>nx7477);
   ix7341 : nor02ii port map ( Y=>nx7340, A0=>nx7727, A1=>nx7481);
   ix7365 : nor02ii port map ( Y=>nx7364, A0=>nx7186, A1=>nx7485);
   ix7395 : nor02ii port map ( Y=>nx7394, A0=>nx7186, A1=>nx7489);
   ix7419 : nor02ii port map ( Y=>nx7418, A0=>nx7186, A1=>nx7493);
   ix7443 : nor02ii port map ( Y=>nx7442, A0=>nx7186, A1=>nx7497);
   ix7467 : nor02ii port map ( Y=>nx7466, A0=>nx7186, A1=>nx7501);
   ix7491 : nor02ii port map ( Y=>nx7490, A0=>nx7186, A1=>nx7505);
   i8_r14_lat_q_13 : latch port map ( Q=>DecompressedData2(223), D=>nx7504, 
      CLK=>nx7731);
   ix7505 : nor02ii port map ( Y=>nx7504, A0=>nx7186, A1=>nx7509);
   ix1193 : nor02ii port map ( Y=>nx1192, A0=>nx7451, A1=>nx1188);
   ix1177 : nand02 port map ( Y=>nx1176, A0=>nx5209, A1=>nx7857);
   ix5210 : nand04 port map ( Y=>nx5209, A0=>nx5121, A1=>nx3895, A2=>nx7439, 
      A3=>nx4665);
   ix1187 : nand02 port map ( Y=>nx1186, A0=>nx5212, A1=>nx5215);
   ix5213 : nand03 port map ( Y=>nx5212, A0=>nx4665, A1=>nx5121, A2=>nx7423
   );
   ix5216 : nor03_2x port map ( Y=>nx5215, A0=>nx1174, A1=>nx7431, A2=>
      nx7407);
   ix1175 : nor02_2x port map ( Y=>nx1174, A0=>nx520, A1=>nx4673);
   ix1207 : nor02ii port map ( Y=>nx1206, A0=>nx7451, A1=>nx1202);
   ix1221 : nor02ii port map ( Y=>nx1220, A0=>nx7451, A1=>nx1216);
   ix1235 : nor02ii port map ( Y=>nx1234, A0=>nx7451, A1=>nx1230);
   ix1249 : nor02ii port map ( Y=>nx1248, A0=>nx7451, A1=>nx1244);
   ix1263 : nor02ii port map ( Y=>nx1262, A0=>nx7451, A1=>nx1258);
   ix1277 : nor02ii port map ( Y=>nx1276, A0=>nx7451, A1=>nx1272);
   ix1291 : nor02ii port map ( Y=>nx1290, A0=>nx1176, A1=>nx1286);
   ix1305 : nor02ii port map ( Y=>nx1304, A0=>nx1176, A1=>nx1300);
   ix1319 : nor02ii port map ( Y=>nx1318, A0=>nx1176, A1=>nx1314);
   ix1333 : nor02ii port map ( Y=>nx1332, A0=>nx1176, A1=>nx1328);
   ix1347 : nor02ii port map ( Y=>nx1346, A0=>nx1176, A1=>nx1342);
   ix1361 : nor02ii port map ( Y=>nx1360, A0=>nx1176, A1=>nx1356);
   ix1375 : nor02ii port map ( Y=>nx1374, A0=>nx1176, A1=>nx1370);
   ix1389 : inv02 port map ( Y=>nx1388, A=>nx5259);
   ix5260 : nor03_2x port map ( Y=>nx5259, A0=>nx1386, A1=>nx7431, A2=>
      nx7409);
   ix1387 : nor02ii port map ( Y=>nx1386, A0=>nx4011, A1=>nx5263);
   ix5264 : nor03_2x port map ( Y=>nx5263, A0=>nx3940, A1=>nx4126, A2=>nx520
   );
   ix1395 : nand02 port map ( Y=>nx1394, A0=>nx5266, A1=>nx5259);
   ix5267 : nand02 port map ( Y=>nx5266, A0=>nx5263, A1=>nx7425);
   ix2087 : nor04 port map ( Y=>nx2086, A0=>nx4532, A1=>nx7839, A2=>nx7447, 
      A3=>nx7409);
   ix2081 : nand02 port map ( Y=>nx2080, A0=>nx5303, A1=>nx7869);
   ix5304 : nand03 port map ( Y=>nx5303, A0=>nx5305, A1=>nx7529, A2=>nx2072
   );
   ix5306 : nor02_2x port map ( Y=>nx5305, A0=>nx4309, A1=>nx4317);
   ix2069 : nor03_2x port map ( Y=>nx2068, A0=>nx7845, A1=>nx4283, A2=>
      nx7839);
   ix2073 : nor02_2x port map ( Y=>nx2072, A0=>nx4318, A1=>i7_counterout2_2
   );
   ix2135 : nor04 port map ( Y=>nx2134, A0=>nx4547, A1=>nx7839, A2=>nx7447, 
      A3=>nx7409);
   ix2161 : nor04 port map ( Y=>nx2160, A0=>nx4553, A1=>nx7841, A2=>nx7447, 
      A3=>nx7409);
   ix2187 : nor04 port map ( Y=>nx2186, A0=>nx4558, A1=>nx7841, A2=>nx7447, 
      A3=>nx7409);
   ix2213 : nor04 port map ( Y=>nx2212, A0=>nx4565, A1=>nx7841, A2=>nx7447, 
      A3=>nx7409);
   ix2239 : nor04 port map ( Y=>nx2238, A0=>nx4570, A1=>nx7841, A2=>nx7447, 
      A3=>nx7411);
   ix2265 : nor04 port map ( Y=>nx2264, A0=>nx4577, A1=>nx7841, A2=>nx7449, 
      A3=>nx7411);
   ix2291 : nor04 port map ( Y=>nx2290, A0=>nx4582, A1=>nx7841, A2=>nx7449, 
      A3=>nx7411);
   ix2321 : nand02 port map ( Y=>nx2320, A0=>nx5331, A1=>nx7869);
   ix5332 : nand03 port map ( Y=>nx5331, A0=>nx5333, A1=>nx7529, A2=>nx2072
   );
   ix5334 : nor02_2x port map ( Y=>nx5333, A0=>i7_counterout2_0, A1=>nx4317
   );
   i7_r27_lat_q_5 : latch port map ( Q=>DecompressedData1(13), D=>nx7553, 
      CLK=>nx7571);
   i7_r27_lat_q_6 : latch port map ( Q=>DecompressedData1(14), D=>nx7559, 
      CLK=>nx7571);
   i7_r27_lat_q_7 : latch port map ( Q=>DecompressedData1(15), D=>nx7565, 
      CLK=>nx7571);
   ix2495 : nand02 port map ( Y=>nx2494, A0=>nx5347, A1=>nx7869);
   ix5348 : nand03 port map ( Y=>nx5347, A0=>nx5349, A1=>nx7529, A2=>nx2072
   );
   ix5350 : nor02_2x port map ( Y=>nx5349, A0=>nx4309, A1=>i7_counterout2_1
   );
   ix2709 : nand02 port map ( Y=>nx2708, A0=>nx5362, A1=>nx7869);
   ix5363 : nand03 port map ( Y=>nx5362, A0=>nx7837, A1=>nx7529, A2=>nx2072
   );
   i7_r25_lat_q_5 : latch port map ( Q=>DecompressedData1(29), D=>nx7553, 
      CLK=>nx7583);
   i7_r25_lat_q_6 : latch port map ( Q=>DecompressedData1(30), D=>nx7559, 
      CLK=>nx7583);
   i7_r25_lat_q_7 : latch port map ( Q=>DecompressedData1(31), D=>nx7565, 
      CLK=>nx7583);
   ix2889 : nand02 port map ( Y=>nx2888, A0=>nx5375, A1=>nx7869);
   ix5376 : nand03 port map ( Y=>nx5375, A0=>nx5305, A1=>nx7529, A2=>nx2880
   );
   ix2881 : nor02_2x port map ( Y=>nx2880, A0=>i7_counterout2_3, A1=>nx4239
   );
   ix3099 : nand02 port map ( Y=>nx3098, A0=>nx5389, A1=>nx7869);
   ix5390 : nand03 port map ( Y=>nx5389, A0=>nx5333, A1=>nx7529, A2=>nx2880
   );
   i7_r23_lat_q_5 : latch port map ( Q=>DecompressedData1(45), D=>nx7553, 
      CLK=>nx7595);
   i7_r23_lat_q_6 : latch port map ( Q=>DecompressedData1(46), D=>nx7559, 
      CLK=>nx7595);
   i7_r23_lat_q_7 : latch port map ( Q=>DecompressedData1(47), D=>nx7565, 
      CLK=>nx7595);
   ix3273 : nand02 port map ( Y=>nx3272, A0=>nx5403, A1=>nx7869);
   ix5404 : nand03 port map ( Y=>nx5403, A0=>nx5349, A1=>nx7529, A2=>nx2880
   );
   ix3487 : nand02 port map ( Y=>nx3486, A0=>nx5415, A1=>nx7871);
   ix5416 : nand03 port map ( Y=>nx5415, A0=>nx7837, A1=>nx7531, A2=>nx2880
   );
   i7_r21_lat_q_5 : latch port map ( Q=>DecompressedData1(61), D=>nx7553, 
      CLK=>nx7607);
   i7_r21_lat_q_6 : latch port map ( Q=>DecompressedData1(62), D=>nx7559, 
      CLK=>nx7607);
   i7_r21_lat_q_7 : latch port map ( Q=>DecompressedData1(63), D=>nx7565, 
      CLK=>nx7607);
   ix3669 : nand02 port map ( Y=>nx3668, A0=>nx5427, A1=>nx7871);
   ix5428 : nand03 port map ( Y=>nx5427, A0=>nx5305, A1=>nx7531, A2=>nx3660
   );
   ix3661 : nor02_2x port map ( Y=>nx3660, A0=>i7_counterout2_3, A1=>
      i7_counterout2_2);
   ix3887 : nand02 port map ( Y=>nx3886, A0=>nx5441, A1=>nx7871);
   ix5442 : nand03 port map ( Y=>nx5441, A0=>nx5333, A1=>nx7531, A2=>nx3660
   );
   i7_r19_lat_q_5 : latch port map ( Q=>DecompressedData1(77), D=>nx7553, 
      CLK=>nx7619);
   i7_r19_lat_q_6 : latch port map ( Q=>DecompressedData1(78), D=>nx7559, 
      CLK=>nx7619);
   i7_r19_lat_q_7 : latch port map ( Q=>DecompressedData1(79), D=>nx7565, 
      CLK=>nx7619);
   ix4061 : nand02 port map ( Y=>nx4060, A0=>nx5454, A1=>nx7871);
   ix5455 : nand03 port map ( Y=>nx5454, A0=>nx5349, A1=>nx7531, A2=>nx3660
   );
   ix4271 : nand02 port map ( Y=>nx4270, A0=>nx5467, A1=>nx7871);
   ix5468 : nand03 port map ( Y=>nx5467, A0=>nx7837, A1=>nx7531, A2=>nx3660
   );
   i7_r17_lat_q_5 : latch port map ( Q=>DecompressedData1(93), D=>nx7553, 
      CLK=>nx7631);
   i7_r17_lat_q_6 : latch port map ( Q=>DecompressedData1(94), D=>nx7559, 
      CLK=>nx7631);
   i7_r17_lat_q_7 : latch port map ( Q=>DecompressedData1(95), D=>nx7565, 
      CLK=>nx7631);
   ix4455 : nand02 port map ( Y=>nx4454, A0=>nx5481, A1=>nx7871);
   ix5482 : nand03 port map ( Y=>nx5481, A0=>nx5305, A1=>nx7635, A2=>nx4446
   );
   ix4447 : nor02_2x port map ( Y=>nx4446, A0=>nx4318, A1=>nx4239);
   ix4665 : nand02 port map ( Y=>nx4664, A0=>nx5497, A1=>nx7871);
   ix5498 : nand03 port map ( Y=>nx5497, A0=>nx5333, A1=>nx7635, A2=>nx4446
   );
   i7_r15_lat_q_5 : latch port map ( Q=>DecompressedData1(109), D=>nx7553, 
      CLK=>nx7651);
   i7_r15_lat_q_6 : latch port map ( Q=>DecompressedData1(110), D=>nx7559, 
      CLK=>nx7651);
   i7_r15_lat_q_7 : latch port map ( Q=>DecompressedData1(111), D=>nx7565, 
      CLK=>nx7651);
   ix4839 : nand02 port map ( Y=>nx4838, A0=>nx5509, A1=>nx7873);
   ix5510 : nand03 port map ( Y=>nx5509, A0=>nx5349, A1=>nx7635, A2=>nx4446
   );
   ix5049 : nand02 port map ( Y=>nx5048, A0=>nx5522, A1=>nx7873);
   ix5523 : nand03 port map ( Y=>nx5522, A0=>nx7837, A1=>nx7635, A2=>nx4446
   );
   i7_r13_lat_q_5 : latch port map ( Q=>DecompressedData1(125), D=>nx7555, 
      CLK=>nx7663);
   i7_r13_lat_q_6 : latch port map ( Q=>DecompressedData1(126), D=>nx7561, 
      CLK=>nx7663);
   i7_r13_lat_q_7 : latch port map ( Q=>DecompressedData1(127), D=>nx7567, 
      CLK=>nx7663);
   ix5229 : nand02 port map ( Y=>nx5228, A0=>nx5535, A1=>nx7873);
   ix5536 : nand03 port map ( Y=>nx5535, A0=>nx5305, A1=>nx7635, A2=>nx5220
   );
   ix5221 : nor02_2x port map ( Y=>nx5220, A0=>nx4318, A1=>i7_counterout2_2
   );
   ix5447 : nand02 port map ( Y=>nx5446, A0=>nx5549, A1=>nx7873);
   ix5550 : nand03 port map ( Y=>nx5549, A0=>nx5333, A1=>nx7635, A2=>nx5220
   );
   i7_r11_lat_q_5 : latch port map ( Q=>DecompressedData1(141), D=>nx7555, 
      CLK=>nx7675);
   i7_r11_lat_q_6 : latch port map ( Q=>DecompressedData1(142), D=>nx7561, 
      CLK=>nx7675);
   i7_r11_lat_q_7 : latch port map ( Q=>DecompressedData1(143), D=>nx7567, 
      CLK=>nx7675);
   ix5621 : nand02 port map ( Y=>nx5620, A0=>nx5562, A1=>nx7873);
   ix5563 : nand03 port map ( Y=>nx5562, A0=>nx5349, A1=>nx7637, A2=>nx5220
   );
   ix5831 : nand02 port map ( Y=>nx5830, A0=>nx5576, A1=>nx7873);
   ix5577 : nand03 port map ( Y=>nx5576, A0=>nx7837, A1=>nx7637, A2=>nx5220
   );
   i7_r9_lat_q_5 : latch port map ( Q=>DecompressedData1(157), D=>nx7555, 
      CLK=>nx7687);
   i7_r9_lat_q_6 : latch port map ( Q=>DecompressedData1(158), D=>nx7561, 
      CLK=>nx7687);
   i7_r9_lat_q_7 : latch port map ( Q=>DecompressedData1(159), D=>nx7567, 
      CLK=>nx7687);
   ix6011 : nand02 port map ( Y=>nx6010, A0=>nx5589, A1=>nx7873);
   ix5590 : nand03 port map ( Y=>nx5589, A0=>nx5305, A1=>nx7637, A2=>nx6002
   );
   ix6003 : nor02_2x port map ( Y=>nx6002, A0=>i7_counterout2_3, A1=>nx4239
   );
   ix6221 : nand02 port map ( Y=>nx6220, A0=>nx5603, A1=>nx7875);
   ix5604 : nand03 port map ( Y=>nx5603, A0=>nx5333, A1=>nx7637, A2=>nx6002
   );
   i7_r7_lat_q_5 : latch port map ( Q=>DecompressedData1(173), D=>nx7555, 
      CLK=>nx7699);
   i7_r7_lat_q_6 : latch port map ( Q=>DecompressedData1(174), D=>nx7561, 
      CLK=>nx7699);
   i7_r7_lat_q_7 : latch port map ( Q=>DecompressedData1(175), D=>nx7567, 
      CLK=>nx7699);
   ix6395 : nand02 port map ( Y=>nx6394, A0=>nx5615, A1=>nx7875);
   ix5616 : nand03 port map ( Y=>nx5615, A0=>nx5349, A1=>nx7637, A2=>nx6002
   );
   ix6605 : nand02 port map ( Y=>nx6604, A0=>nx5628, A1=>nx7875);
   ix5629 : nand03 port map ( Y=>nx5628, A0=>nx4293, A1=>nx7637, A2=>nx6002
   );
   i7_r5_lat_q_5 : latch port map ( Q=>DecompressedData1(189), D=>nx7555, 
      CLK=>nx7711);
   i7_r5_lat_q_6 : latch port map ( Q=>DecompressedData1(190), D=>nx7561, 
      CLK=>nx7711);
   i7_r5_lat_q_7 : latch port map ( Q=>DecompressedData1(191), D=>nx7567, 
      CLK=>nx7711);
   ix6787 : nand02 port map ( Y=>nx6786, A0=>nx5643, A1=>nx7875);
   ix5644 : nand03 port map ( Y=>nx5643, A0=>nx5305, A1=>nx7639, A2=>nx6778
   );
   ix6779 : nor02_2x port map ( Y=>nx6778, A0=>i7_counterout2_3, A1=>
      i7_counterout2_2);
   ix6997 : nand02 port map ( Y=>nx6996, A0=>nx5659, A1=>nx7875);
   ix5660 : nand03 port map ( Y=>nx5659, A0=>nx5333, A1=>nx7639, A2=>nx6778
   );
   i7_r3_lat_q_5 : latch port map ( Q=>DecompressedData1(205), D=>nx7555, 
      CLK=>nx7723);
   i7_r3_lat_q_6 : latch port map ( Q=>DecompressedData1(206), D=>nx7561, 
      CLK=>nx7723);
   i7_r3_lat_q_7 : latch port map ( Q=>DecompressedData1(207), D=>nx7567, 
      CLK=>nx7723);
   ix7171 : nand02 port map ( Y=>nx7170, A0=>nx5671, A1=>nx7875);
   ix5672 : nand03 port map ( Y=>nx5671, A0=>nx5349, A1=>nx7639, A2=>nx6778
   );
   ix7381 : nand02 port map ( Y=>nx7380, A0=>nx5684, A1=>nx7875);
   ix5685 : nand03 port map ( Y=>nx5684, A0=>nx4293, A1=>nx7639, A2=>nx6778
   );
   i7_r1_lat_q_5 : latch port map ( Q=>DecompressedData1(221), D=>nx7555, 
      CLK=>nx7735);
   i7_r1_lat_q_6 : latch port map ( Q=>DecompressedData1(222), D=>nx7561, 
      CLK=>nx7735);
   i7_r1_lat_q_7 : latch port map ( Q=>DecompressedData1(223), D=>nx7567, 
      CLK=>nx7735);
   ix2133 : mux21 port map ( Y=>DecompressedData(0), A0=>nx5695, A1=>nx5697, 
      S0=>CNNIMGLOAD);
   ix2159 : mux21 port map ( Y=>DecompressedData(1), A0=>nx5700, A1=>nx5703, 
      S0=>CNNIMGLOAD);
   ix2185 : mux21 port map ( Y=>DecompressedData(2), A0=>nx5707, A1=>nx5709, 
      S0=>CNNIMGLOAD);
   ix2211 : mux21 port map ( Y=>DecompressedData(3), A0=>nx5712, A1=>nx5715, 
      S0=>CNNIMGLOAD);
   ix2237 : mux21 port map ( Y=>DecompressedData(4), A0=>nx5719, A1=>nx5721, 
      S0=>CNNIMGLOAD);
   ix2263 : mux21 port map ( Y=>DecompressedData(5), A0=>nx5724, A1=>nx5727, 
      S0=>CNNIMGLOAD);
   ix2289 : mux21 port map ( Y=>DecompressedData(6), A0=>nx5731, A1=>nx5733, 
      S0=>CNNIMGLOAD);
   ix2315 : mux21 port map ( Y=>DecompressedData(7), A0=>nx5736, A1=>nx5739, 
      S0=>CNNIMGLOAD);
   ix2345 : mux21 port map ( Y=>DecompressedData(8), A0=>nx5743, A1=>nx5745, 
      S0=>CNNIMGLOAD);
   ix2369 : mux21 port map ( Y=>DecompressedData(9), A0=>nx5748, A1=>nx5751, 
      S0=>CNNIMGLOAD);
   ix2393 : mux21 port map ( Y=>DecompressedData(10), A0=>nx5755, A1=>nx5757, 
      S0=>CNNIMGLOAD);
   ix2417 : mux21 port map ( Y=>DecompressedData(11), A0=>nx5760, A1=>nx5763, 
      S0=>CNNIMGLOAD);
   ix2441 : mux21 port map ( Y=>DecompressedData(12), A0=>nx5767, A1=>nx5769, 
      S0=>CNNIMGLOAD);
   ix2465 : nand02 port map ( Y=>DecompressedData(13), A0=>nx5772, A1=>
      nx5775);
   ix5773 : nand02 port map ( Y=>nx5772, A0=>nx7743, A1=>
      DecompressedData1(13));
   ix5776 : nand02 port map ( Y=>nx5775, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(15));
   ix2477 : nand02 port map ( Y=>DecompressedData(14), A0=>nx5779, A1=>
      nx5775);
   ix5780 : nand02 port map ( Y=>nx5779, A0=>nx7743, A1=>
      DecompressedData1(14));
   ix2489 : nand02 port map ( Y=>DecompressedData(15), A0=>nx5782, A1=>
      nx5775);
   ix5783 : nand02 port map ( Y=>nx5782, A0=>nx7743, A1=>
      DecompressedData1(15));
   ix2535 : mux21 port map ( Y=>DecompressedData(16), A0=>nx5785, A1=>nx5787, 
      S0=>CNNIMGLOAD);
   ix2559 : mux21 port map ( Y=>DecompressedData(17), A0=>nx5791, A1=>nx5793, 
      S0=>CNNIMGLOAD);
   ix2583 : mux21 port map ( Y=>DecompressedData(18), A0=>nx5796, A1=>nx5799, 
      S0=>CNNIMGLOAD);
   ix2607 : mux21 port map ( Y=>DecompressedData(19), A0=>nx5803, A1=>nx5805, 
      S0=>CNNIMGLOAD);
   ix2631 : mux21 port map ( Y=>DecompressedData(20), A0=>nx5808, A1=>nx5811, 
      S0=>CNNIMGLOAD);
   ix2655 : mux21 port map ( Y=>DecompressedData(21), A0=>nx5815, A1=>nx5817, 
      S0=>CNNIMGLOAD);
   ix2679 : mux21 port map ( Y=>DecompressedData(22), A0=>nx5820, A1=>nx5823, 
      S0=>CNNIMGLOAD);
   ix2703 : mux21 port map ( Y=>DecompressedData(23), A0=>nx5827, A1=>nx5829, 
      S0=>CNNIMGLOAD);
   ix2733 : mux21 port map ( Y=>DecompressedData(24), A0=>nx5833, A1=>nx5835, 
      S0=>CNNIMGLOAD);
   ix2757 : mux21 port map ( Y=>DecompressedData(25), A0=>nx5838, A1=>nx5841, 
      S0=>CNNIMGLOAD);
   ix2781 : mux21 port map ( Y=>DecompressedData(26), A0=>nx5845, A1=>nx5847, 
      S0=>CNNIMGLOAD);
   ix2805 : mux21 port map ( Y=>DecompressedData(27), A0=>nx5850, A1=>nx5853, 
      S0=>CNNIMGLOAD);
   ix2829 : mux21 port map ( Y=>DecompressedData(28), A0=>nx5857, A1=>nx5859, 
      S0=>CNNIMGLOAD);
   ix2853 : nand02 port map ( Y=>DecompressedData(29), A0=>nx5862, A1=>
      nx5865);
   ix5863 : nand02 port map ( Y=>nx5862, A0=>nx7743, A1=>
      DecompressedData1(29));
   ix5866 : nand02 port map ( Y=>nx5865, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(31));
   ix2865 : nand02 port map ( Y=>DecompressedData(30), A0=>nx5869, A1=>
      nx5865);
   ix5870 : nand02 port map ( Y=>nx5869, A0=>nx7743, A1=>
      DecompressedData1(30));
   ix2877 : nand02 port map ( Y=>DecompressedData(31), A0=>nx5872, A1=>
      nx5865);
   ix5873 : nand02 port map ( Y=>nx5872, A0=>nx7743, A1=>
      DecompressedData1(31));
   ix2925 : mux21 port map ( Y=>DecompressedData(32), A0=>nx5875, A1=>nx5877, 
      S0=>CNNIMGLOAD);
   ix2949 : mux21 port map ( Y=>DecompressedData(33), A0=>nx5881, A1=>nx5883, 
      S0=>CNNIMGLOAD);
   ix2973 : mux21 port map ( Y=>DecompressedData(34), A0=>nx5886, A1=>nx5889, 
      S0=>CNNIMGLOAD);
   ix2997 : mux21 port map ( Y=>DecompressedData(35), A0=>nx5893, A1=>nx5895, 
      S0=>CNNIMGLOAD);
   ix3021 : mux21 port map ( Y=>DecompressedData(36), A0=>nx5898, A1=>nx5901, 
      S0=>CNNIMGLOAD);
   ix3045 : mux21 port map ( Y=>DecompressedData(37), A0=>nx5905, A1=>nx5907, 
      S0=>CNNIMGLOAD);
   ix3069 : mux21 port map ( Y=>DecompressedData(38), A0=>nx5910, A1=>nx5913, 
      S0=>CNNIMGLOAD);
   ix3093 : mux21 port map ( Y=>DecompressedData(39), A0=>nx5917, A1=>nx5919, 
      S0=>CNNIMGLOAD);
   ix3123 : mux21 port map ( Y=>DecompressedData(40), A0=>nx5922, A1=>nx5925, 
      S0=>CNNIMGLOAD);
   ix3147 : mux21 port map ( Y=>DecompressedData(41), A0=>nx5929, A1=>nx5931, 
      S0=>CNNIMGLOAD);
   ix3171 : mux21 port map ( Y=>DecompressedData(42), A0=>nx5934, A1=>nx5937, 
      S0=>CNNIMGLOAD);
   ix3195 : mux21 port map ( Y=>DecompressedData(43), A0=>nx5941, A1=>nx5943, 
      S0=>CNNIMGLOAD);
   ix3219 : mux21 port map ( Y=>DecompressedData(44), A0=>nx5946, A1=>nx5949, 
      S0=>CNNIMGLOAD);
   ix3243 : nand02 port map ( Y=>DecompressedData(45), A0=>nx5953, A1=>
      nx5955);
   ix5954 : nand02 port map ( Y=>nx5953, A0=>nx7745, A1=>
      DecompressedData1(45));
   ix5956 : nand02 port map ( Y=>nx5955, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(47));
   ix3255 : nand02 port map ( Y=>DecompressedData(46), A0=>nx5958, A1=>
      nx5955);
   ix5959 : nand02 port map ( Y=>nx5958, A0=>nx7745, A1=>
      DecompressedData1(46));
   ix3267 : nand02 port map ( Y=>DecompressedData(47), A0=>nx5961, A1=>
      nx5955);
   ix5962 : nand02 port map ( Y=>nx5961, A0=>nx7745, A1=>
      DecompressedData1(47));
   ix3313 : mux21 port map ( Y=>DecompressedData(48), A0=>nx5965, A1=>nx5967, 
      S0=>CNNIMGLOAD);
   ix3337 : mux21 port map ( Y=>DecompressedData(49), A0=>nx5970, A1=>nx5973, 
      S0=>CNNIMGLOAD);
   ix3361 : mux21 port map ( Y=>DecompressedData(50), A0=>nx5977, A1=>nx5979, 
      S0=>CNNIMGLOAD);
   ix3385 : mux21 port map ( Y=>DecompressedData(51), A0=>nx5982, A1=>nx5985, 
      S0=>CNNIMGLOAD);
   ix3409 : mux21 port map ( Y=>DecompressedData(52), A0=>nx5989, A1=>nx5991, 
      S0=>CNNIMGLOAD);
   ix3433 : mux21 port map ( Y=>DecompressedData(53), A0=>nx5994, A1=>nx5997, 
      S0=>CNNIMGLOAD);
   ix3457 : mux21 port map ( Y=>DecompressedData(54), A0=>nx6001, A1=>nx6003, 
      S0=>CNNIMGLOAD);
   ix3481 : mux21 port map ( Y=>DecompressedData(55), A0=>nx6007, A1=>nx6009, 
      S0=>CNNIMGLOAD);
   ix3511 : mux21 port map ( Y=>DecompressedData(56), A0=>nx6013, A1=>nx6015, 
      S0=>CNNIMGLOAD);
   ix3535 : mux21 port map ( Y=>DecompressedData(57), A0=>nx6018, A1=>nx6021, 
      S0=>CNNIMGLOAD);
   ix3559 : mux21 port map ( Y=>DecompressedData(58), A0=>nx6025, A1=>nx6027, 
      S0=>CNNIMGLOAD);
   ix3583 : mux21 port map ( Y=>DecompressedData(59), A0=>nx6031, A1=>nx6033, 
      S0=>CNNIMGLOAD);
   ix3607 : mux21 port map ( Y=>DecompressedData(60), A0=>nx6037, A1=>nx6039, 
      S0=>CNNIMGLOAD);
   ix3631 : nand02 port map ( Y=>DecompressedData(61), A0=>nx6042, A1=>
      nx6045);
   ix6043 : nand02 port map ( Y=>nx6042, A0=>nx7745, A1=>
      DecompressedData1(61));
   ix6046 : nand02 port map ( Y=>nx6045, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(63));
   ix3643 : nand02 port map ( Y=>DecompressedData(62), A0=>nx6049, A1=>
      nx6045);
   ix6050 : nand02 port map ( Y=>nx6049, A0=>nx7745, A1=>
      DecompressedData1(62));
   ix3655 : nand02 port map ( Y=>DecompressedData(63), A0=>nx6052, A1=>
      nx6045);
   ix6053 : nand02 port map ( Y=>nx6052, A0=>nx7745, A1=>
      DecompressedData1(63));
   ix3713 : mux21 port map ( Y=>DecompressedData(64), A0=>nx6055, A1=>nx6057, 
      S0=>CNNIMGLOAD);
   ix3737 : mux21 port map ( Y=>DecompressedData(65), A0=>nx6061, A1=>nx6063, 
      S0=>CNNIMGLOAD);
   ix3761 : mux21 port map ( Y=>DecompressedData(66), A0=>nx6066, A1=>nx6069, 
      S0=>CNNIMGLOAD);
   ix3785 : mux21 port map ( Y=>DecompressedData(67), A0=>nx6073, A1=>nx6075, 
      S0=>CNNIMGLOAD);
   ix3809 : mux21 port map ( Y=>DecompressedData(68), A0=>nx6078, A1=>nx6081, 
      S0=>CNNIMGLOAD);
   ix3833 : mux21 port map ( Y=>DecompressedData(69), A0=>nx6085, A1=>nx6087, 
      S0=>CNNIMGLOAD);
   ix3857 : mux21 port map ( Y=>DecompressedData(70), A0=>nx6090, A1=>nx6093, 
      S0=>CNNIMGLOAD);
   ix3881 : mux21 port map ( Y=>DecompressedData(71), A0=>nx6097, A1=>nx6099, 
      S0=>CNNIMGLOAD);
   ix3911 : mux21 port map ( Y=>DecompressedData(72), A0=>nx6102, A1=>nx6105, 
      S0=>CNNIMGLOAD);
   ix3935 : mux21 port map ( Y=>DecompressedData(73), A0=>nx6109, A1=>nx6111, 
      S0=>CNNIMGLOAD);
   ix3959 : mux21 port map ( Y=>DecompressedData(74), A0=>nx6114, A1=>nx6117, 
      S0=>CNNIMGLOAD);
   ix3983 : mux21 port map ( Y=>DecompressedData(75), A0=>nx6121, A1=>nx6123, 
      S0=>CNNIMGLOAD);
   ix4007 : mux21 port map ( Y=>DecompressedData(76), A0=>nx6126, A1=>nx6129, 
      S0=>CNNIMGLOAD);
   ix4031 : nand02 port map ( Y=>DecompressedData(77), A0=>nx6133, A1=>
      nx6135);
   ix6134 : nand02 port map ( Y=>nx6133, A0=>nx7745, A1=>
      DecompressedData1(77));
   ix6136 : nand02 port map ( Y=>nx6135, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(79));
   ix4043 : nand02 port map ( Y=>DecompressedData(78), A0=>nx6138, A1=>
      nx6135);
   ix6139 : nand02 port map ( Y=>nx6138, A0=>nx7747, A1=>
      DecompressedData1(78));
   ix4055 : nand02 port map ( Y=>DecompressedData(79), A0=>nx6141, A1=>
      nx6135);
   ix6142 : nand02 port map ( Y=>nx6141, A0=>nx7747, A1=>
      DecompressedData1(79));
   ix4097 : mux21 port map ( Y=>DecompressedData(80), A0=>nx6145, A1=>nx6147, 
      S0=>CNNIMGLOAD);
   ix4121 : mux21 port map ( Y=>DecompressedData(81), A0=>nx6150, A1=>nx6153, 
      S0=>CNNIMGLOAD);
   ix4145 : mux21 port map ( Y=>DecompressedData(82), A0=>nx6157, A1=>nx6159, 
      S0=>CNNIMGLOAD);
   ix4169 : mux21 port map ( Y=>DecompressedData(83), A0=>nx6162, A1=>nx6165, 
      S0=>CNNIMGLOAD);
   ix4193 : mux21 port map ( Y=>DecompressedData(84), A0=>nx6169, A1=>nx6171, 
      S0=>CNNIMGLOAD);
   ix4217 : mux21 port map ( Y=>DecompressedData(85), A0=>nx6174, A1=>nx6177, 
      S0=>CNNIMGLOAD);
   ix4241 : mux21 port map ( Y=>DecompressedData(86), A0=>nx6181, A1=>nx6183, 
      S0=>CNNIMGLOAD);
   ix4265 : mux21 port map ( Y=>DecompressedData(87), A0=>nx6186, A1=>nx6189, 
      S0=>CNNIMGLOAD);
   ix4295 : mux21 port map ( Y=>DecompressedData(88), A0=>nx6193, A1=>nx6195, 
      S0=>CNNIMGLOAD);
   ix4319 : mux21 port map ( Y=>DecompressedData(89), A0=>nx6198, A1=>nx6201, 
      S0=>CNNIMGLOAD);
   ix4343 : mux21 port map ( Y=>DecompressedData(90), A0=>nx6205, A1=>nx6207, 
      S0=>CNNIMGLOAD);
   ix4367 : mux21 port map ( Y=>DecompressedData(91), A0=>nx6210, A1=>nx6213, 
      S0=>CNNIMGLOAD);
   ix4391 : mux21 port map ( Y=>DecompressedData(92), A0=>nx6217, A1=>nx6219, 
      S0=>CNNIMGLOAD);
   ix4415 : nand02 port map ( Y=>DecompressedData(93), A0=>nx6223, A1=>
      nx6225);
   ix6224 : nand02 port map ( Y=>nx6223, A0=>nx7747, A1=>
      DecompressedData1(93));
   ix6226 : nand02 port map ( Y=>nx6225, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(95));
   ix4427 : nand02 port map ( Y=>DecompressedData(94), A0=>nx6228, A1=>
      nx6225);
   ix6229 : nand02 port map ( Y=>nx6228, A0=>nx7747, A1=>
      DecompressedData1(94));
   ix4439 : nand02 port map ( Y=>DecompressedData(95), A0=>nx6231, A1=>
      nx6225);
   ix6232 : nand02 port map ( Y=>nx6231, A0=>nx7747, A1=>
      DecompressedData1(95));
   ix4491 : mux21 port map ( Y=>DecompressedData(96), A0=>nx6235, A1=>nx6237, 
      S0=>CNNIMGLOAD);
   ix4515 : mux21 port map ( Y=>DecompressedData(97), A0=>nx6240, A1=>nx6243, 
      S0=>CNNIMGLOAD);
   ix4539 : mux21 port map ( Y=>DecompressedData(98), A0=>nx6247, A1=>nx6249, 
      S0=>CNNIMGLOAD);
   ix4563 : mux21 port map ( Y=>DecompressedData(99), A0=>nx6252, A1=>nx6255, 
      S0=>CNNIMGLOAD);
   ix4587 : mux21 port map ( Y=>DecompressedData(100), A0=>nx6259, A1=>
      nx6261, S0=>CNNIMGLOAD);
   ix4611 : mux21 port map ( Y=>DecompressedData(101), A0=>nx6264, A1=>
      nx6267, S0=>CNNIMGLOAD);
   ix4635 : mux21 port map ( Y=>DecompressedData(102), A0=>nx6271, A1=>
      nx6273, S0=>CNNIMGLOAD);
   ix4659 : mux21 port map ( Y=>DecompressedData(103), A0=>nx6276, A1=>
      nx6279, S0=>CNNIMGLOAD);
   ix4689 : mux21 port map ( Y=>DecompressedData(104), A0=>nx6283, A1=>
      nx6285, S0=>CNNIMGLOAD);
   ix4713 : mux21 port map ( Y=>DecompressedData(105), A0=>nx6288, A1=>
      nx6291, S0=>CNNIMGLOAD);
   ix4737 : mux21 port map ( Y=>DecompressedData(106), A0=>nx6295, A1=>
      nx6297, S0=>CNNIMGLOAD);
   ix4761 : mux21 port map ( Y=>DecompressedData(107), A0=>nx6300, A1=>
      nx6303, S0=>CNNIMGLOAD);
   ix4785 : mux21 port map ( Y=>DecompressedData(108), A0=>nx6307, A1=>
      nx6309, S0=>CNNIMGLOAD);
   ix4809 : nand02 port map ( Y=>DecompressedData(109), A0=>nx6312, A1=>
      nx6315);
   ix6313 : nand02 port map ( Y=>nx6312, A0=>nx7747, A1=>
      DecompressedData1(109));
   ix6316 : nand02 port map ( Y=>nx6315, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(111));
   ix4821 : nand02 port map ( Y=>DecompressedData(110), A0=>nx6319, A1=>
      nx6315);
   ix6320 : nand02 port map ( Y=>nx6319, A0=>nx7747, A1=>
      DecompressedData1(110));
   ix4833 : nand02 port map ( Y=>DecompressedData(111), A0=>nx6322, A1=>
      nx6315);
   ix6323 : nand02 port map ( Y=>nx6322, A0=>nx7749, A1=>
      DecompressedData1(111));
   ix4875 : mux21 port map ( Y=>DecompressedData(112), A0=>nx6325, A1=>
      nx6327, S0=>CNNIMGLOAD);
   ix4899 : mux21 port map ( Y=>DecompressedData(113), A0=>nx6331, A1=>
      nx6333, S0=>CNNIMGLOAD);
   ix4923 : mux21 port map ( Y=>DecompressedData(114), A0=>nx6336, A1=>
      nx6339, S0=>CNNIMGLOAD);
   ix4947 : mux21 port map ( Y=>DecompressedData(115), A0=>nx6343, A1=>
      nx6345, S0=>CNNIMGLOAD);
   ix4971 : mux21 port map ( Y=>DecompressedData(116), A0=>nx6348, A1=>
      nx6350, S0=>CNNIMGLOAD);
   ix4995 : mux21 port map ( Y=>DecompressedData(117), A0=>nx6353, A1=>
      nx6355, S0=>CNNIMGLOAD);
   ix5019 : mux21 port map ( Y=>DecompressedData(118), A0=>nx6358, A1=>
      nx6360, S0=>CNNIMGLOAD);
   ix5043 : mux21 port map ( Y=>DecompressedData(119), A0=>nx6363, A1=>
      nx6365, S0=>CNNIMGLOAD);
   ix5073 : mux21 port map ( Y=>DecompressedData(120), A0=>nx6368, A1=>
      nx6370, S0=>CNNIMGLOAD);
   ix5097 : mux21 port map ( Y=>DecompressedData(121), A0=>nx6373, A1=>
      nx6375, S0=>CNNIMGLOAD);
   ix5121 : mux21 port map ( Y=>DecompressedData(122), A0=>nx6379, A1=>
      nx6381, S0=>CNNIMGLOAD);
   ix5145 : mux21 port map ( Y=>DecompressedData(123), A0=>nx6384, A1=>
      nx6387, S0=>CNNIMGLOAD);
   ix5169 : mux21 port map ( Y=>DecompressedData(124), A0=>nx6391, A1=>
      nx6393, S0=>CNNIMGLOAD);
   ix5193 : nand02 port map ( Y=>DecompressedData(125), A0=>nx6397, A1=>
      nx6399);
   ix6398 : nand02 port map ( Y=>nx6397, A0=>nx7749, A1=>
      DecompressedData1(125));
   ix6400 : nand02 port map ( Y=>nx6399, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(127));
   ix5205 : nand02 port map ( Y=>DecompressedData(126), A0=>nx6402, A1=>
      nx6399);
   ix6403 : nand02 port map ( Y=>nx6402, A0=>nx7749, A1=>
      DecompressedData1(126));
   ix5217 : nand02 port map ( Y=>DecompressedData(127), A0=>nx6405, A1=>
      nx6399);
   ix6406 : nand02 port map ( Y=>nx6405, A0=>nx7749, A1=>
      DecompressedData1(127));
   ix5273 : mux21 port map ( Y=>DecompressedData(128), A0=>nx6409, A1=>
      nx6411, S0=>CNNIMGLOAD);
   ix5297 : mux21 port map ( Y=>DecompressedData(129), A0=>nx6415, A1=>
      nx6417, S0=>CNNIMGLOAD);
   ix5321 : mux21 port map ( Y=>DecompressedData(130), A0=>nx6421, A1=>
      nx6423, S0=>CNNIMGLOAD);
   ix5345 : mux21 port map ( Y=>DecompressedData(131), A0=>nx6426, A1=>
      nx6429, S0=>CNNIMGLOAD);
   ix5369 : mux21 port map ( Y=>DecompressedData(132), A0=>nx6433, A1=>
      nx6435, S0=>CNNIMGLOAD);
   ix5393 : mux21 port map ( Y=>DecompressedData(133), A0=>nx6438, A1=>
      nx6441, S0=>CNNIMGLOAD);
   ix5417 : mux21 port map ( Y=>DecompressedData(134), A0=>nx6445, A1=>
      nx6447, S0=>CNNIMGLOAD);
   ix5441 : mux21 port map ( Y=>DecompressedData(135), A0=>nx6450, A1=>
      nx6453, S0=>CNNIMGLOAD);
   ix5471 : mux21 port map ( Y=>DecompressedData(136), A0=>nx6457, A1=>
      nx6459, S0=>CNNIMGLOAD);
   ix5495 : mux21 port map ( Y=>DecompressedData(137), A0=>nx6462, A1=>
      nx6465, S0=>CNNIMGLOAD);
   ix5519 : mux21 port map ( Y=>DecompressedData(138), A0=>nx6469, A1=>
      nx6471, S0=>CNNIMGLOAD);
   ix5543 : mux21 port map ( Y=>DecompressedData(139), A0=>nx6474, A1=>
      nx6477, S0=>CNNIMGLOAD);
   ix5567 : mux21 port map ( Y=>DecompressedData(140), A0=>nx6481, A1=>
      nx6483, S0=>CNNIMGLOAD);
   ix5591 : nand02 port map ( Y=>DecompressedData(141), A0=>nx6486, A1=>
      nx6489);
   ix6487 : nand02 port map ( Y=>nx6486, A0=>nx7749, A1=>
      DecompressedData1(141));
   ix6490 : nand02 port map ( Y=>nx6489, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(143));
   ix5603 : nand02 port map ( Y=>DecompressedData(142), A0=>nx6493, A1=>
      nx6489);
   ix6494 : nand02 port map ( Y=>nx6493, A0=>nx7749, A1=>
      DecompressedData1(142));
   ix5615 : nand02 port map ( Y=>DecompressedData(143), A0=>nx6496, A1=>
      nx6489);
   ix6497 : nand02 port map ( Y=>nx6496, A0=>nx7749, A1=>
      DecompressedData1(143));
   ix5657 : mux21 port map ( Y=>DecompressedData(144), A0=>nx6499, A1=>
      nx6501, S0=>CNNIMGLOAD);
   ix5681 : mux21 port map ( Y=>DecompressedData(145), A0=>nx6505, A1=>
      nx6507, S0=>CNNIMGLOAD);
   ix5705 : mux21 port map ( Y=>DecompressedData(146), A0=>nx6510, A1=>
      nx6513, S0=>CNNIMGLOAD);
   ix5729 : mux21 port map ( Y=>DecompressedData(147), A0=>nx6517, A1=>
      nx6519, S0=>CNNIMGLOAD);
   ix5753 : mux21 port map ( Y=>DecompressedData(148), A0=>nx6522, A1=>
      nx6525, S0=>CNNIMGLOAD);
   ix5777 : mux21 port map ( Y=>DecompressedData(149), A0=>nx6529, A1=>
      nx6531, S0=>CNNIMGLOAD);
   ix5801 : mux21 port map ( Y=>DecompressedData(150), A0=>nx6534, A1=>
      nx6537, S0=>CNNIMGLOAD);
   ix5825 : mux21 port map ( Y=>DecompressedData(151), A0=>nx6541, A1=>
      nx6543, S0=>CNNIMGLOAD);
   ix5855 : mux21 port map ( Y=>DecompressedData(152), A0=>nx6546, A1=>
      nx6549, S0=>CNNIMGLOAD);
   ix5879 : mux21 port map ( Y=>DecompressedData(153), A0=>nx6553, A1=>
      nx6555, S0=>CNNIMGLOAD);
   ix5903 : mux21 port map ( Y=>DecompressedData(154), A0=>nx6558, A1=>
      nx6561, S0=>CNNIMGLOAD);
   ix5927 : mux21 port map ( Y=>DecompressedData(155), A0=>nx6565, A1=>
      nx6567, S0=>CNNIMGLOAD);
   ix5951 : mux21 port map ( Y=>DecompressedData(156), A0=>nx6570, A1=>
      nx6573, S0=>CNNIMGLOAD);
   ix5975 : nand02 port map ( Y=>DecompressedData(157), A0=>nx6577, A1=>
      nx6579);
   ix6578 : nand02 port map ( Y=>nx6577, A0=>nx7751, A1=>
      DecompressedData1(157));
   ix6580 : nand02 port map ( Y=>nx6579, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(159));
   ix5987 : nand02 port map ( Y=>DecompressedData(158), A0=>nx6582, A1=>
      nx6579);
   ix6583 : nand02 port map ( Y=>nx6582, A0=>nx7751, A1=>
      DecompressedData1(158));
   ix5999 : nand02 port map ( Y=>DecompressedData(159), A0=>nx6585, A1=>
      nx6579);
   ix6586 : nand02 port map ( Y=>nx6585, A0=>nx7751, A1=>
      DecompressedData1(159));
   ix6047 : mux21 port map ( Y=>DecompressedData(160), A0=>nx6589, A1=>
      nx6591, S0=>CNNIMGLOAD);
   ix6071 : mux21 port map ( Y=>DecompressedData(161), A0=>nx6594, A1=>
      nx6597, S0=>CNNIMGLOAD);
   ix6095 : mux21 port map ( Y=>DecompressedData(162), A0=>nx6601, A1=>
      nx6603, S0=>CNNIMGLOAD);
   ix6119 : mux21 port map ( Y=>DecompressedData(163), A0=>nx6607, A1=>
      nx6609, S0=>CNNIMGLOAD);
   ix6143 : mux21 port map ( Y=>DecompressedData(164), A0=>nx6612, A1=>
      nx6615, S0=>CNNIMGLOAD);
   ix6167 : mux21 port map ( Y=>DecompressedData(165), A0=>nx6619, A1=>
      nx6621, S0=>CNNIMGLOAD);
   ix6191 : mux21 port map ( Y=>DecompressedData(166), A0=>nx6624, A1=>
      nx6627, S0=>CNNIMGLOAD);
   ix6215 : mux21 port map ( Y=>DecompressedData(167), A0=>nx6631, A1=>
      nx6633, S0=>CNNIMGLOAD);
   ix6245 : mux21 port map ( Y=>DecompressedData(168), A0=>nx6636, A1=>
      nx6639, S0=>CNNIMGLOAD);
   ix6269 : mux21 port map ( Y=>DecompressedData(169), A0=>nx6643, A1=>
      nx6645, S0=>CNNIMGLOAD);
   ix6293 : mux21 port map ( Y=>DecompressedData(170), A0=>nx6648, A1=>
      nx6651, S0=>CNNIMGLOAD);
   ix6317 : mux21 port map ( Y=>DecompressedData(171), A0=>nx6655, A1=>
      nx6657, S0=>CNNIMGLOAD);
   ix6341 : mux21 port map ( Y=>DecompressedData(172), A0=>nx6660, A1=>
      nx6663, S0=>CNNIMGLOAD);
   ix6365 : nand02 port map ( Y=>DecompressedData(173), A0=>nx6667, A1=>
      nx6669);
   ix6668 : nand02 port map ( Y=>nx6667, A0=>nx7751, A1=>
      DecompressedData1(173));
   ix6670 : nand02 port map ( Y=>nx6669, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(175));
   ix6377 : nand02 port map ( Y=>DecompressedData(174), A0=>nx6672, A1=>
      nx6669);
   ix6673 : nand02 port map ( Y=>nx6672, A0=>nx7751, A1=>
      DecompressedData1(174));
   ix6389 : nand02 port map ( Y=>DecompressedData(175), A0=>nx6675, A1=>
      nx6669);
   ix6676 : nand02 port map ( Y=>nx6675, A0=>nx7751, A1=>
      DecompressedData1(175));
   ix6431 : mux21 port map ( Y=>DecompressedData(176), A0=>nx6679, A1=>
      nx6681, S0=>CNNIMGLOAD);
   ix6455 : mux21 port map ( Y=>DecompressedData(177), A0=>nx6684, A1=>
      nx6687, S0=>CNNIMGLOAD);
   ix6479 : mux21 port map ( Y=>DecompressedData(178), A0=>nx6691, A1=>
      nx6693, S0=>CNNIMGLOAD);
   ix6503 : mux21 port map ( Y=>DecompressedData(179), A0=>nx6696, A1=>
      nx6699, S0=>CNNIMGLOAD);
   ix6527 : mux21 port map ( Y=>DecompressedData(180), A0=>nx6703, A1=>
      nx6705, S0=>CNNIMGLOAD);
   ix6551 : mux21 port map ( Y=>DecompressedData(181), A0=>nx6708, A1=>
      nx6711, S0=>CNNIMGLOAD);
   ix6575 : mux21 port map ( Y=>DecompressedData(182), A0=>nx6715, A1=>
      nx6717, S0=>CNNIMGLOAD);
   ix6599 : mux21 port map ( Y=>DecompressedData(183), A0=>nx6720, A1=>
      nx6723, S0=>CNNIMGLOAD);
   ix6629 : mux21 port map ( Y=>DecompressedData(184), A0=>nx6727, A1=>
      nx6729, S0=>CNNIMGLOAD);
   ix6653 : mux21 port map ( Y=>DecompressedData(185), A0=>nx6732, A1=>
      nx6734, S0=>CNNIMGLOAD);
   ix6677 : mux21 port map ( Y=>DecompressedData(186), A0=>nx6737, A1=>
      nx6739, S0=>CNNIMGLOAD);
   ix6701 : mux21 port map ( Y=>DecompressedData(187), A0=>nx6742, A1=>
      nx6744, S0=>CNNIMGLOAD);
   ix6725 : mux21 port map ( Y=>DecompressedData(188), A0=>nx6747, A1=>
      nx6749, S0=>CNNIMGLOAD);
   ix6749 : nand02 port map ( Y=>DecompressedData(189), A0=>nx6752, A1=>
      nx6754);
   ix6753 : nand02 port map ( Y=>nx6752, A0=>nx7751, A1=>
      DecompressedData1(189));
   ix6755 : nand02 port map ( Y=>nx6754, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(191));
   ix6761 : nand02 port map ( Y=>DecompressedData(190), A0=>nx6757, A1=>
      nx6754);
   ix6758 : nand02 port map ( Y=>nx6757, A0=>nx7753, A1=>
      DecompressedData1(190));
   ix6773 : nand02 port map ( Y=>DecompressedData(191), A0=>nx6761, A1=>
      nx6754);
   ix6762 : nand02 port map ( Y=>nx6761, A0=>nx7753, A1=>
      DecompressedData1(191));
   ix6823 : mux21 port map ( Y=>DecompressedData(192), A0=>nx6764, A1=>
      nx6766, S0=>CNNIMGLOAD);
   ix6847 : mux21 port map ( Y=>DecompressedData(193), A0=>nx6769, A1=>
      nx6771, S0=>CNNIMGLOAD);
   ix6871 : mux21 port map ( Y=>DecompressedData(194), A0=>nx6775, A1=>
      nx6777, S0=>CNNIMGLOAD);
   ix6895 : mux21 port map ( Y=>DecompressedData(195), A0=>nx6781, A1=>
      nx6783, S0=>CNNIMGLOAD);
   ix6919 : mux21 port map ( Y=>DecompressedData(196), A0=>nx6787, A1=>
      nx6789, S0=>CNNIMGLOAD);
   ix6943 : mux21 port map ( Y=>DecompressedData(197), A0=>nx6792, A1=>
      nx6794, S0=>CNNIMGLOAD);
   ix6967 : mux21 port map ( Y=>DecompressedData(198), A0=>nx6797, A1=>
      nx6799, S0=>CNNIMGLOAD);
   ix6991 : mux21 port map ( Y=>DecompressedData(199), A0=>nx6803, A1=>
      nx6805, S0=>CNNIMGLOAD);
   ix7021 : mux21 port map ( Y=>DecompressedData(200), A0=>nx6809, A1=>
      nx6811, S0=>CNNIMGLOAD);
   ix7045 : mux21 port map ( Y=>DecompressedData(201), A0=>nx6815, A1=>
      nx6817, S0=>CNNIMGLOAD);
   ix7069 : mux21 port map ( Y=>DecompressedData(202), A0=>nx6821, A1=>
      nx6823, S0=>CNNIMGLOAD);
   ix7093 : mux21 port map ( Y=>DecompressedData(203), A0=>nx6826, A1=>
      nx6828, S0=>CNNIMGLOAD);
   ix7117 : mux21 port map ( Y=>DecompressedData(204), A0=>nx6831, A1=>
      nx6833, S0=>CNNIMGLOAD);
   ix7141 : nand02 port map ( Y=>DecompressedData(205), A0=>nx6837, A1=>
      nx6839);
   ix6838 : nand02 port map ( Y=>nx6837, A0=>nx7753, A1=>
      DecompressedData1(205));
   ix6840 : nand02 port map ( Y=>nx6839, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(207));
   ix7153 : nand02 port map ( Y=>DecompressedData(206), A0=>nx6842, A1=>
      nx6839);
   ix6843 : nand02 port map ( Y=>nx6842, A0=>nx7753, A1=>
      DecompressedData1(206));
   ix7165 : nand02 port map ( Y=>DecompressedData(207), A0=>nx6845, A1=>
      nx6839);
   ix6846 : nand02 port map ( Y=>nx6845, A0=>nx7753, A1=>
      DecompressedData1(207));
   ix7207 : mux21 port map ( Y=>DecompressedData(208), A0=>nx6849, A1=>
      nx6851, S0=>CNNIMGLOAD);
   ix7231 : mux21 port map ( Y=>DecompressedData(209), A0=>nx6854, A1=>
      nx6857, S0=>CNNIMGLOAD);
   ix7255 : mux21 port map ( Y=>DecompressedData(210), A0=>nx6861, A1=>
      nx6863, S0=>CNNIMGLOAD);
   ix7279 : mux21 port map ( Y=>DecompressedData(211), A0=>nx6866, A1=>
      nx6869, S0=>CNNIMGLOAD);
   ix7303 : mux21 port map ( Y=>DecompressedData(212), A0=>nx6873, A1=>
      nx6875, S0=>CNNIMGLOAD);
   ix7327 : mux21 port map ( Y=>DecompressedData(213), A0=>nx6878, A1=>
      nx6881, S0=>CNNIMGLOAD);
   ix7351 : mux21 port map ( Y=>DecompressedData(214), A0=>nx6885, A1=>
      nx6887, S0=>CNNIMGLOAD);
   ix7375 : mux21 port map ( Y=>DecompressedData(215), A0=>nx6890, A1=>
      nx6893, S0=>CNNIMGLOAD);
   ix7405 : mux21 port map ( Y=>DecompressedData(216), A0=>nx6897, A1=>
      nx6899, S0=>CNNIMGLOAD);
   ix7429 : mux21 port map ( Y=>DecompressedData(217), A0=>nx6902, A1=>
      nx6905, S0=>CNNIMGLOAD);
   ix7453 : mux21 port map ( Y=>DecompressedData(218), A0=>nx6909, A1=>
      nx6911, S0=>CNNIMGLOAD);
   ix7477 : mux21 port map ( Y=>DecompressedData(219), A0=>nx6914, A1=>
      nx6917, S0=>CNNIMGLOAD);
   ix7501 : mux21 port map ( Y=>DecompressedData(220), A0=>nx6921, A1=>
      nx6923, S0=>CNNIMGLOAD);
   ix7525 : nand02 port map ( Y=>DecompressedData(221), A0=>nx6926, A1=>
      nx6929);
   ix6927 : nand02 port map ( Y=>nx6926, A0=>nx7753, A1=>
      DecompressedData1(221));
   ix6930 : nand02 port map ( Y=>nx6929, A0=>CNNIMGLOAD, A1=>
      DecompressedData2(223));
   ix7537 : nand02 port map ( Y=>DecompressedData(222), A0=>nx6933, A1=>
      nx6929);
   ix6934 : nand02 port map ( Y=>nx6933, A0=>nx7753, A1=>
      DecompressedData1(222));
   ix7549 : nand02 port map ( Y=>DecompressedData(223), A0=>nx6936, A1=>
      nx6929);
   ix6937 : nand02 port map ( Y=>nx6936, A0=>nx7755, A1=>
      DecompressedData1(223));
   ix1201 : nor02_2x port map ( Y=>DecompressedData(224), A0=>nx7755, A1=>
      nx6939);
   ix1215 : nor02_2x port map ( Y=>DecompressedData(225), A0=>nx7755, A1=>
      nx6943);
   ix1229 : nor02_2x port map ( Y=>DecompressedData(226), A0=>nx7755, A1=>
      nx6946);
   ix1243 : nor02_2x port map ( Y=>DecompressedData(227), A0=>nx7755, A1=>
      nx6949);
   ix1257 : nor02_2x port map ( Y=>DecompressedData(228), A0=>nx7755, A1=>
      nx6953);
   ix1271 : nor02_2x port map ( Y=>DecompressedData(229), A0=>nx7755, A1=>
      nx6957);
   ix1285 : nor02_2x port map ( Y=>DecompressedData(230), A0=>nx7757, A1=>
      nx6960);
   ix1299 : nor02_2x port map ( Y=>DecompressedData(231), A0=>nx7757, A1=>
      nx6963);
   ix1313 : nor02_2x port map ( Y=>DecompressedData(232), A0=>nx7757, A1=>
      nx6967);
   ix1327 : nor02_2x port map ( Y=>DecompressedData(233), A0=>nx7757, A1=>
      nx6970);
   ix1341 : nor02_2x port map ( Y=>DecompressedData(234), A0=>nx7757, A1=>
      nx6973);
   ix1355 : nor02_2x port map ( Y=>DecompressedData(235), A0=>nx7757, A1=>
      nx6977);
   ix1369 : nor02_2x port map ( Y=>DecompressedData(236), A0=>nx7757, A1=>
      nx6981);
   ix1383 : nor02_2x port map ( Y=>DecompressedData(239), A0=>nx7759, A1=>
      nx6984);
   ix1407 : nor02_2x port map ( Y=>DecompressedData(240), A0=>nx7759, A1=>
      nx6987);
   ix1419 : nor02_2x port map ( Y=>DecompressedData(241), A0=>nx7759, A1=>
      nx6991);
   ix1431 : nor02_2x port map ( Y=>DecompressedData(242), A0=>nx7759, A1=>
      nx6995);
   ix1443 : nor02_2x port map ( Y=>DecompressedData(243), A0=>nx7759, A1=>
      nx6999);
   ix1455 : nor02_2x port map ( Y=>DecompressedData(244), A0=>nx7759, A1=>
      nx7002);
   ix1467 : nor02_2x port map ( Y=>DecompressedData(245), A0=>nx7759, A1=>
      nx7005);
   ix1479 : nor02_2x port map ( Y=>DecompressedData(246), A0=>nx7761, A1=>
      nx7009);
   ix1491 : nor02_2x port map ( Y=>DecompressedData(247), A0=>nx7761, A1=>
      nx7013);
   ix1503 : nor02_2x port map ( Y=>DecompressedData(248), A0=>nx7761, A1=>
      nx7016);
   ix1515 : nor02_2x port map ( Y=>DecompressedData(249), A0=>nx7761, A1=>
      nx7019);
   ix1527 : nor02_2x port map ( Y=>DecompressedData(250), A0=>nx7761, A1=>
      nx7023);
   ix1539 : nor02_2x port map ( Y=>DecompressedData(251), A0=>nx7761, A1=>
      nx7026);
   ix1551 : nor02_2x port map ( Y=>DecompressedData(252), A0=>nx7761, A1=>
      nx7029);
   ix1563 : nor02_2x port map ( Y=>DecompressedData(255), A0=>nx7763, A1=>
      nx7033);
   ix7038 : inv01 port map ( Y=>nx7037, A=>OuterAddress(0));
   i5_aa_reg_Q : dff port map ( Q=>i5_FAEN, QB=>OPEN, D=>nx1616, CLK=>CLK);
   ix1617 : nor02ii port map ( Y=>nx1616, A0=>nx7045, A1=>nx1614);
   ix7046 : nor02_2x port map ( Y=>nx7045, A0=>nx1606, A1=>nx1604);
   ix1607 : nor02_2x port map ( Y=>nx1606, A0=>nx7957, A1=>nx7048);
   ix7049 : aoi21 port map ( Y=>nx7048, A0=>OuterWrite, A1=>
      ProcessEnable_EXMPLR, B0=>DecompressionDone);
   ix1595 : nand02 port map ( Y=>DecompressionDone, A0=>nx7051, A1=>nx7057);
   i7_reg_readtoRam : dffs_ni port map ( Q=>DecompressionDone1, QB=>nx7051, 
      D=>nx3503, CLK=>CLK, S=>NOT_nx814);
   ix3504 : nor02_2x port map ( Y=>nx3503, A0=>nx7051, A1=>nx814);
   i8_reg_ramWrite : dffs_ni port map ( Q=>DecompressionDone2, QB=>nx7057, D
      =>nx3493, CLK=>CLK, S=>nx558);
   ix3494 : nor02_2x port map ( Y=>nx3493, A0=>nx7057, A1=>nx546);
   ix559 : nand02 port map ( Y=>nx558, A0=>nx546, A1=>nx4011);
   ix1605 : nor03_2x port map ( Y=>nx1604, A0=>nx3563, A1=>nx7063, A2=>
      nx1598);
   ix7064 : inv01 port map ( Y=>nx7063, A=>INCEnable);
   ix1599 : nand03 port map ( Y=>nx1598, A0=>nx7067, A1=>nx7051, A2=>nx7057
   );
   ix7068 : nand02 port map ( Y=>nx7067, A0=>OuterWrite, A1=>
      ProcessEnable_EXMPLR);
   ix1615 : nor02_2x port map ( Y=>nx1614, A0=>Rst, A1=>nx7515);
   i5_MR_reg_dataout_0 : dffr port map ( Q=>i5_MARo_0, QB=>nx7039, D=>nx1634, 
      CLK=>CLK, R=>Rst);
   ix7080 : inv01 port map ( Y=>nx7079, A=>OuterAddress(1));
   i5_MR_reg_dataout_1 : dffr port map ( Q=>i5_MARo_1, QB=>nx7081, D=>nx1660, 
      CLK=>CLK, R=>Rst);
   ix1661 : oai21 port map ( Y=>nx1660, A0=>nx7877, A1=>nx7085, B0=>nx7088);
   ix7086 : xnor2 port map ( Y=>nx7085, A0=>nx1626, A1=>Address(1));
   ix1627 : nand02 port map ( Y=>nx1626, A0=>nx7072, A1=>nx7515);
   ix7089 : oai21 port map ( Y=>nx7088, A0=>nx1670, A1=>nx1668, B0=>nx7877);
   ix1671 : nor02_2x port map ( Y=>nx1670, A0=>nx7079, A1=>nx7889);
   ix1669 : nor02_2x port map ( Y=>nx1668, A0=>nx7081, A1=>nx7521);
   ix1643 : nor02_2x port map ( Y=>nx1642, A0=>nx7095, A1=>nx7907);
   ix7096 : inv01 port map ( Y=>nx7095, A=>ActivateOuterAddress);
   ix7099 : inv01 port map ( Y=>nx7098, A=>OuterAddress(2));
   i5_MR_reg_dataout_2 : dffr port map ( Q=>i5_MARo_2, QB=>nx7100, D=>nx1688, 
      CLK=>CLK, R=>Rst);
   ix1689 : oai21 port map ( Y=>nx1688, A0=>nx7877, A1=>nx7103, B0=>nx7109);
   ix7104 : xnor2 port map ( Y=>nx7103, A0=>nx1682, A1=>Address(2));
   ix1683 : oai21 port map ( Y=>nx1682, A0=>nx7072, A1=>nx7107, B0=>nx7515);
   ix7110 : oai21 port map ( Y=>nx7109, A0=>nx1698, A1=>nx1696, B0=>nx7877);
   ix1699 : nor02_2x port map ( Y=>nx1698, A0=>nx7098, A1=>nx7889);
   ix1697 : nor02_2x port map ( Y=>nx1696, A0=>nx7100, A1=>nx7521);
   ix7116 : inv01 port map ( Y=>nx7115, A=>OuterAddress(3));
   ix1717 : oai21 port map ( Y=>nx1716, A0=>nx7877, A1=>nx7121, B0=>nx7132);
   ix7122 : xnor2 port map ( Y=>nx7121, A0=>nx7123, A1=>nx7129);
   ix7124 : nand02 port map ( Y=>nx7123, A0=>nx1682, A1=>nx1708);
   ix1709 : nand02 port map ( Y=>nx1708, A0=>nx7126, A1=>nx7515);
   i5_MR_reg_dataout_3 : dffr port map ( Q=>i5_MARo_3, QB=>nx7117, D=>nx1716, 
      CLK=>CLK, R=>Rst);
   ix7133 : oai21 port map ( Y=>nx7132, A0=>nx1726, A1=>nx1724, B0=>nx7877);
   ix1727 : nor02_2x port map ( Y=>nx1726, A0=>nx7115, A1=>nx7891);
   ix1725 : nor02_2x port map ( Y=>nx1724, A0=>nx7117, A1=>nx7521);
   ix7138 : inv01 port map ( Y=>nx7137, A=>OuterAddress(4));
   ix1745 : oai21 port map ( Y=>nx1744, A0=>nx7877, A1=>nx7143, B0=>nx7151);
   ix7144 : xnor2 port map ( Y=>nx7143, A0=>nx7145, A1=>nx7148);
   ix7146 : nand03 port map ( Y=>nx7145, A0=>nx1682, A1=>nx1708, A2=>nx1736
   );
   ix1737 : nand02 port map ( Y=>nx1736, A0=>nx7129, A1=>nx7515);
   i5_MR_reg_dataout_4 : dffr port map ( Q=>i5_MARo_4, QB=>nx7139, D=>nx1744, 
      CLK=>CLK, R=>Rst);
   ix7152 : oai21 port map ( Y=>nx7151, A0=>nx1754, A1=>nx1752, B0=>nx7879);
   ix1755 : nor02_2x port map ( Y=>nx1754, A0=>nx7137, A1=>nx7891);
   ix1753 : nor02_2x port map ( Y=>nx1752, A0=>nx7139, A1=>nx7521);
   ix7158 : inv01 port map ( Y=>nx7157, A=>OuterAddress(5));
   ix1773 : oai21 port map ( Y=>nx1772, A0=>nx7879, A1=>nx7163, B0=>nx7173);
   ix7164 : xnor2 port map ( Y=>nx7163, A0=>nx7165, A1=>nx7169);
   ix7166 : nand04 port map ( Y=>nx7165, A0=>nx1682, A1=>nx1708, A2=>nx1736, 
      A3=>nx1764);
   ix1765 : nand02 port map ( Y=>nx1764, A0=>nx7148, A1=>nx7515);
   i5_MR_reg_dataout_5 : dffr port map ( Q=>i5_MARo_5, QB=>nx7159, D=>nx1772, 
      CLK=>CLK, R=>Rst);
   ix7174 : oai21 port map ( Y=>nx7173, A0=>nx1782, A1=>nx1780, B0=>nx7879);
   ix1783 : nor02_2x port map ( Y=>nx1782, A0=>nx7157, A1=>nx7893);
   ix1781 : nor02_2x port map ( Y=>nx1780, A0=>nx7159, A1=>nx7521);
   ix7179 : inv01 port map ( Y=>nx7178, A=>OuterAddress(6));
   i5_MR_reg_dataout_6 : dffr port map ( Q=>i5_MARo_6, QB=>nx7181, D=>nx1800, 
      CLK=>CLK, R=>Rst);
   ix1801 : oai21 port map ( Y=>nx1800, A0=>nx7879, A1=>nx7185, B0=>nx7189);
   ix7186 : xnor2 port map ( Y=>nx7185, A0=>nx7525, A1=>Address(6));
   ix1795 : aoi21 port map ( Y=>nx1794, A0=>nx7169, A1=>nx7517, B0=>nx7165);
   ix7190 : oai21 port map ( Y=>nx7189, A0=>nx1810, A1=>nx1808, B0=>nx7879);
   ix1811 : nor02_2x port map ( Y=>nx1810, A0=>nx7178, A1=>nx7893);
   ix1809 : nor02_2x port map ( Y=>nx1808, A0=>nx7181, A1=>nx7521);
   ix7198 : inv01 port map ( Y=>nx7197, A=>OuterAddress(7));
   ix1829 : oai21 port map ( Y=>nx1828, A0=>nx7879, A1=>nx7202, B0=>nx7214);
   ix7203 : xnor2 port map ( Y=>nx7202, A0=>nx7205, A1=>nx7211);
   ix7206 : nand02 port map ( Y=>nx7205, A0=>nx7525, A1=>nx1820);
   ix1821 : nand02 port map ( Y=>nx1820, A0=>nx7209, A1=>nx7517);
   i5_MR_reg_dataout_7 : dffr port map ( Q=>i5_MARo_7, QB=>nx7199, D=>nx1828, 
      CLK=>CLK, R=>Rst);
   ix7215 : oai21 port map ( Y=>nx7214, A0=>nx1838, A1=>nx1836, B0=>nx7879);
   ix1839 : nor02_2x port map ( Y=>nx1838, A0=>nx7197, A1=>nx7895);
   ix1837 : nor02_2x port map ( Y=>nx1836, A0=>nx7199, A1=>nx7523);
   ix7222 : inv01 port map ( Y=>nx7221, A=>OuterAddress(8));
   ix1857 : oai21 port map ( Y=>nx1856, A0=>nx7881, A1=>nx7226, B0=>nx7236);
   ix7227 : xnor2 port map ( Y=>nx7226, A0=>nx7229, A1=>nx7233);
   ix7230 : nand03 port map ( Y=>nx7229, A0=>nx7525, A1=>nx1820, A2=>nx1848
   );
   ix1849 : nand02 port map ( Y=>nx1848, A0=>nx7211, A1=>nx7517);
   i5_MR_reg_dataout_8 : dffr port map ( Q=>i5_MARo_8, QB=>nx7223, D=>nx1856, 
      CLK=>CLK, R=>Rst);
   ix7237 : oai21 port map ( Y=>nx7236, A0=>nx1866, A1=>nx1864, B0=>nx7881);
   ix1867 : nor02_2x port map ( Y=>nx1866, A0=>nx7221, A1=>nx7895);
   ix1865 : nor02_2x port map ( Y=>nx1864, A0=>nx7223, A1=>nx7523);
   ix7242 : inv01 port map ( Y=>nx7241, A=>OuterAddress(9));
   ix1885 : oai21 port map ( Y=>nx1884, A0=>nx7881, A1=>nx7247, B0=>nx7257);
   ix7248 : xnor2 port map ( Y=>nx7247, A0=>nx7249, A1=>nx7253);
   ix7250 : nand04 port map ( Y=>nx7249, A0=>nx7525, A1=>nx1820, A2=>nx1848, 
      A3=>nx1876);
   ix1877 : nand02 port map ( Y=>nx1876, A0=>nx7233, A1=>nx7517);
   i5_MR_reg_dataout_9 : dffr port map ( Q=>i5_MARo_9, QB=>nx7243, D=>nx1884, 
      CLK=>CLK, R=>Rst);
   ix7258 : oai21 port map ( Y=>nx7257, A0=>nx1894, A1=>nx1892, B0=>nx7881);
   ix1895 : nor02_2x port map ( Y=>nx1894, A0=>nx7241, A1=>nx7895);
   ix1893 : nor02_2x port map ( Y=>nx1892, A0=>nx7243, A1=>nx7523);
   ix7263 : inv01 port map ( Y=>nx7262, A=>OuterAddress(10));
   i5_MR_reg_dataout_10 : dffr port map ( Q=>i5_MARo_10, QB=>nx7265, D=>
      nx1912, CLK=>CLK, R=>Rst);
   ix1913 : oai21 port map ( Y=>nx1912, A0=>nx7881, A1=>nx7269, B0=>nx7272);
   ix7270 : xnor2 port map ( Y=>nx7269, A0=>nx7527, A1=>Address(10));
   ix1907 : aoi21 port map ( Y=>nx1906, A0=>nx7253, A1=>nx7517, B0=>nx7249);
   ix7273 : oai21 port map ( Y=>nx7272, A0=>nx1922, A1=>nx1920, B0=>nx7881);
   ix1923 : nor02_2x port map ( Y=>nx1922, A0=>nx7262, A1=>nx7897);
   ix1921 : nor02_2x port map ( Y=>nx1920, A0=>nx7265, A1=>nx7523);
   ix7278 : inv01 port map ( Y=>nx7277, A=>OuterAddress(11));
   ix1941 : oai21 port map ( Y=>nx1940, A0=>nx7881, A1=>nx7282, B0=>nx7293);
   ix7283 : xnor2 port map ( Y=>nx7282, A0=>nx7284, A1=>nx7289);
   ix7285 : nand02 port map ( Y=>nx7284, A0=>nx7527, A1=>nx1932);
   ix1933 : nand02 port map ( Y=>nx1932, A0=>nx7287, A1=>nx7517);
   i5_MR_reg_dataout_11 : dffr port map ( Q=>i5_MARo_11, QB=>nx7279, D=>
      nx1940, CLK=>CLK, R=>Rst);
   ix7294 : oai21 port map ( Y=>nx7293, A0=>nx1950, A1=>nx1948, B0=>nx7883);
   ix1951 : nor02_2x port map ( Y=>nx1950, A0=>nx7277, A1=>nx7897);
   ix1949 : nor02_2x port map ( Y=>nx1948, A0=>nx7279, A1=>nx7523);
   ix7299 : inv01 port map ( Y=>nx7298, A=>OuterAddress(12));
   ix1969 : oai21 port map ( Y=>nx1968, A0=>nx7883, A1=>nx7305, B0=>nx7313);
   ix7306 : xnor2 port map ( Y=>nx7305, A0=>nx7307, A1=>nx7310);
   ix7308 : nand03 port map ( Y=>nx7307, A0=>nx7527, A1=>nx1932, A2=>nx1960
   );
   ix1961 : nand02 port map ( Y=>nx1960, A0=>nx7289, A1=>nx7517);
   i5_MR_reg_dataout_12 : dffr port map ( Q=>i5_MARo_12, QB=>nx7301, D=>
      nx1968, CLK=>CLK, R=>Rst);
   ix7314 : oai21 port map ( Y=>nx7313, A0=>nx1978, A1=>nx1976, B0=>nx7883);
   ix1979 : nor02_2x port map ( Y=>nx1978, A0=>nx7298, A1=>nx7899);
   ix1977 : nor02_2x port map ( Y=>nx1976, A0=>nx7301, A1=>nx7523);
   ix7320 : inv01 port map ( Y=>nx7319, A=>OuterAddress(13));
   ix1997 : oai21 port map ( Y=>nx1996, A0=>nx7883, A1=>nx7325, B0=>nx7333);
   ix7326 : xnor2 port map ( Y=>nx7325, A0=>nx7327, A1=>nx7330);
   ix7328 : nand04 port map ( Y=>nx7327, A0=>nx7527, A1=>nx1932, A2=>nx1960, 
      A3=>nx1988);
   ix1989 : nand02 port map ( Y=>nx1988, A0=>nx7310, A1=>nx7519);
   i5_MR_reg_dataout_13 : dffr port map ( Q=>i5_MARo_13, QB=>nx7321, D=>
      nx1996, CLK=>CLK, R=>Rst);
   ix7334 : oai21 port map ( Y=>nx7333, A0=>nx2006, A1=>nx2004, B0=>nx7883);
   ix2007 : nor02_2x port map ( Y=>nx2006, A0=>nx7319, A1=>nx7899);
   ix2005 : nor02_2x port map ( Y=>nx2004, A0=>nx7321, A1=>nx1642);
   ix7340 : inv01 port map ( Y=>nx7339, A=>OuterAddress(14));
   i5_MR_reg_dataout_14 : dffr port map ( Q=>i5_MARo_14, QB=>nx7341, D=>
      nx2024, CLK=>CLK, R=>Rst);
   ix2025 : oai21 port map ( Y=>nx2024, A0=>nx7883, A1=>nx7344, B0=>nx7347);
   ix7345 : xnor2 port map ( Y=>nx7344, A0=>nx2018, A1=>Address(14));
   ix2019 : aoi21 port map ( Y=>nx2018, A0=>nx7330, A1=>nx7519, B0=>nx7327);
   ix7348 : oai21 port map ( Y=>nx7347, A0=>nx2034, A1=>nx2032, B0=>nx7883);
   ix2035 : nor02_2x port map ( Y=>nx2034, A0=>nx7339, A1=>nx7899);
   ix2033 : nor02_2x port map ( Y=>nx2032, A0=>nx7341, A1=>nx1642);
   ix7355 : inv01 port map ( Y=>nx7354, A=>OuterAddress(15));
   ix2053 : oai21 port map ( Y=>nx2052, A0=>nx7885, A1=>nx7359, B0=>nx7370);
   ix7360 : xnor2 port map ( Y=>nx7359, A0=>nx7361, A1=>nx7367);
   ix7362 : nand02 port map ( Y=>nx7361, A0=>nx2018, A1=>nx2044);
   ix2045 : nand02 port map ( Y=>nx2044, A0=>nx7365, A1=>nx7519);
   i5_MR_reg_dataout_15 : dffr port map ( Q=>i5_MARo_15, QB=>nx7356, D=>
      nx2052, CLK=>CLK, R=>Rst);
   ix7371 : oai21 port map ( Y=>nx7370, A0=>nx2062, A1=>nx2060, B0=>nx7885);
   ix2063 : nor02_2x port map ( Y=>nx2062, A0=>nx7354, A1=>nx7901);
   ix2061 : nor02_2x port map ( Y=>nx2060, A0=>nx7356, A1=>nx1642);
   ix7551 : nor02_2x port map ( Y=>readenable, A0=>nx7377, A1=>nx3563);
   ix7378 : inv01 port map ( Y=>nx7377, A=>OuterRead);
   ix1167 : nand02 port map ( Y=>EnableReadingFromCPU, A0=>nx7381, A1=>
      nx7383);
   ix7382 : nand03 port map ( Y=>nx7381, A0=>nx7392, A1=>nx7763, A2=>nx7907
   );
   ix7384 : nand03 port map ( Y=>nx7383, A0=>nx7397, A1=>CNNIMGLOAD, A2=>
      nx7907);
   ix7389 : inv02 port map ( Y=>nx7390, A=>nx4203);
   ix7391 : inv02 port map ( Y=>nx7392, A=>nx4203);
   ix7393 : inv02 port map ( Y=>nx7395, A=>nx4083);
   ix7396 : inv02 port map ( Y=>nx7397, A=>nx4083);
   ix7400 : inv04 port map ( Y=>nx7401, A=>nx7399);
   ix7402 : inv04 port map ( Y=>nx7403, A=>nx9396);
   ix7404 : inv04 port map ( Y=>nx7405, A=>nx9396);
   ix7406 : inv04 port map ( Y=>nx7407, A=>nx9396);
   ix7408 : inv04 port map ( Y=>nx7409, A=>nx9396);
   ix7410 : inv04 port map ( Y=>nx7411, A=>nx9396);
   ix7412 : inv02 port map ( Y=>nx7413, A=>nx7771);
   ix7414 : inv02 port map ( Y=>nx7415, A=>nx7771);
   ix7416 : inv01 port map ( Y=>nx7417, A=>nx370);
   ix7418 : inv02 port map ( Y=>nx7419, A=>nx7417);
   ix7420 : inv02 port map ( Y=>nx7421, A=>nx7417);
   ix7422 : inv02 port map ( Y=>nx7423, A=>nx7417);
   ix7424 : inv02 port map ( Y=>nx7425, A=>nx7417);
   ix7426 : buf02 port map ( Y=>nx7427, A=>nx374);
   ix7428 : buf02 port map ( Y=>nx7429, A=>nx374);
   ix7430 : buf02 port map ( Y=>nx7431, A=>nx374);
   ix7434 : inv02 port map ( Y=>nx7435, A=>nx7433);
   ix7436 : inv02 port map ( Y=>nx7437, A=>nx7433);
   ix7438 : inv02 port map ( Y=>nx7439, A=>nx7433);
   ix7440 : inv02 port map ( Y=>nx7441, A=>nx4217);
   ix7442 : inv02 port map ( Y=>nx7443, A=>nx4217);
   ix7444 : inv02 port map ( Y=>nx7445, A=>nx4217);
   ix7446 : inv02 port map ( Y=>nx7447, A=>nx4301);
   ix7448 : inv02 port map ( Y=>nx7449, A=>nx4301);
   ix7450 : nand02 port map ( Y=>nx7451, A0=>nx5209, A1=>nx7857);
   ix7454 : nor02_2x port map ( Y=>nx7455, A0=>nx4532, A1=>nx7789);
   ix7456 : nor02_2x port map ( Y=>nx7457, A0=>nx4532, A1=>nx7789);
   ix7458 : nor02_2x port map ( Y=>nx7459, A0=>nx4547, A1=>nx7789);
   ix7460 : nor02_2x port map ( Y=>nx7461, A0=>nx4547, A1=>nx7789);
   ix7462 : nor02_2x port map ( Y=>nx7463, A0=>nx4553, A1=>nx7789);
   ix7464 : nor02_2x port map ( Y=>nx7465, A0=>nx4553, A1=>nx7791);
   ix7466 : nor02_2x port map ( Y=>nx7467, A0=>nx4558, A1=>nx7791);
   ix7468 : nor02_2x port map ( Y=>nx7469, A0=>nx4558, A1=>nx7791);
   ix7470 : nor02_2x port map ( Y=>nx7471, A0=>nx4565, A1=>nx7791);
   ix7472 : nor02_2x port map ( Y=>nx7473, A0=>nx4565, A1=>nx7791);
   ix7474 : nor02_2x port map ( Y=>nx7475, A0=>nx4570, A1=>nx7791);
   ix7476 : nor02_2x port map ( Y=>nx7477, A0=>nx4570, A1=>nx7791);
   ix7478 : nor02_2x port map ( Y=>nx7479, A0=>nx4577, A1=>nx7793);
   ix7480 : nor02_2x port map ( Y=>nx7481, A0=>nx4577, A1=>nx7793);
   ix7482 : nor02_2x port map ( Y=>nx7483, A0=>nx4582, A1=>nx7793);
   ix7484 : nor02_2x port map ( Y=>nx7485, A0=>nx4582, A1=>nx7793);
   ix7486 : nor02_2x port map ( Y=>nx7487, A0=>nx4511, A1=>nx7793);
   ix7488 : nor02_2x port map ( Y=>nx7489, A0=>nx4511, A1=>nx7793);
   ix7490 : nor02_2x port map ( Y=>nx7491, A0=>nx4592, A1=>nx7793);
   ix7492 : nor02_2x port map ( Y=>nx7493, A0=>nx4592, A1=>nx7795);
   ix7494 : nor02_2x port map ( Y=>nx7495, A0=>nx4397, A1=>nx7795);
   ix7496 : nor02_2x port map ( Y=>nx7497, A0=>nx4397, A1=>nx7795);
   ix7498 : nor02_2x port map ( Y=>nx7499, A0=>nx4377, A1=>nx7795);
   ix7500 : nor02_2x port map ( Y=>nx7501, A0=>nx4377, A1=>nx7795);
   ix7502 : nor02_2x port map ( Y=>nx7503, A0=>nx4381, A1=>nx7795);
   ix7504 : nor02_2x port map ( Y=>nx7505, A0=>nx4381, A1=>nx7795);
   ix7506 : nor02_2x port map ( Y=>nx7507, A0=>nx4460, A1=>nx7797);
   ix7508 : nor02_2x port map ( Y=>nx7509, A0=>nx4460, A1=>nx7797);
   ix7510 : inv02 port map ( Y=>nx7511, A=>nx5259);
   ix7514 : inv02 port map ( Y=>nx7515, A=>nx7885);
   ix7516 : inv02 port map ( Y=>nx7517, A=>nx7885);
   ix7518 : inv02 port map ( Y=>nx7519, A=>nx7885);
   ix7520 : nor02_2x port map ( Y=>nx7521, A0=>nx7095, A1=>nx7909);
   ix7522 : nor02_2x port map ( Y=>nx7523, A0=>nx7095, A1=>nx7909);
   ix7524 : buf02 port map ( Y=>nx7525, A=>nx1794);
   ix7526 : buf02 port map ( Y=>nx7527, A=>nx1906);
   ix7528 : buf02 port map ( Y=>nx7529, A=>nx2068);
   ix7530 : buf02 port map ( Y=>nx7531, A=>nx2068);
   ix7536 : nand02 port map ( Y=>nx7537, A0=>nx4522, A1=>nx7857);
   ix7538 : inv01 port map ( Y=>nx7539, A=>nx2118);
   ix7540 : inv01 port map ( Y=>nx7541, A=>nx7539);
   ix7550 : inv01 port map ( Y=>nx7551, A=>nx2238);
   ix7552 : inv02 port map ( Y=>nx7553, A=>nx7551);
   ix7554 : inv02 port map ( Y=>nx7555, A=>nx7551);
   ix7556 : inv01 port map ( Y=>nx7557, A=>nx2264);
   ix7558 : inv02 port map ( Y=>nx7559, A=>nx7557);
   ix7560 : inv02 port map ( Y=>nx7561, A=>nx7557);
   ix7562 : inv01 port map ( Y=>nx7563, A=>nx2290);
   ix7564 : inv02 port map ( Y=>nx7565, A=>nx7563);
   ix7566 : inv02 port map ( Y=>nx7567, A=>nx7563);
   ix7568 : inv01 port map ( Y=>nx7569, A=>nx2320);
   ix7570 : inv01 port map ( Y=>nx7571, A=>nx7569);
   ix7574 : nand02 port map ( Y=>nx7575, A0=>nx4613, A1=>nx7857);
   ix7576 : inv01 port map ( Y=>nx7577, A=>nx2520);
   ix7578 : inv01 port map ( Y=>nx7579, A=>nx7577);
   ix7580 : inv01 port map ( Y=>nx7581, A=>nx2708);
   ix7582 : inv01 port map ( Y=>nx7583, A=>nx7581);
   ix7586 : nand02 port map ( Y=>nx7587, A0=>nx4663, A1=>nx7857);
   ix7588 : inv01 port map ( Y=>nx7589, A=>nx2910);
   ix7590 : inv01 port map ( Y=>nx7591, A=>nx7589);
   ix7592 : inv01 port map ( Y=>nx7593, A=>nx3098);
   ix7594 : inv01 port map ( Y=>nx7595, A=>nx7593);
   ix7598 : nand02 port map ( Y=>nx7599, A0=>nx4711, A1=>nx7857);
   ix7600 : inv01 port map ( Y=>nx7601, A=>nx3298);
   ix7602 : inv01 port map ( Y=>nx7603, A=>nx7601);
   ix7604 : inv01 port map ( Y=>nx7605, A=>nx3486);
   ix7606 : inv01 port map ( Y=>nx7607, A=>nx7605);
   ix7610 : nand02 port map ( Y=>nx7611, A0=>nx4757, A1=>nx7857);
   ix7612 : inv01 port map ( Y=>nx7613, A=>nx3698);
   ix7614 : inv01 port map ( Y=>nx7615, A=>nx7613);
   ix7616 : inv01 port map ( Y=>nx7617, A=>nx3886);
   ix7618 : inv01 port map ( Y=>nx7619, A=>nx7617);
   ix7622 : nand02 port map ( Y=>nx7623, A0=>nx4804, A1=>nx7859);
   ix7624 : inv01 port map ( Y=>nx7625, A=>nx4082);
   ix7626 : inv01 port map ( Y=>nx7627, A=>nx7625);
   ix7628 : inv01 port map ( Y=>nx7629, A=>nx4270);
   ix7630 : inv01 port map ( Y=>nx7631, A=>nx7629);
   ix7634 : inv01 port map ( Y=>nx7635, A=>nx7633);
   ix7636 : inv01 port map ( Y=>nx7637, A=>nx7633);
   ix7638 : inv01 port map ( Y=>nx7639, A=>nx7633);
   ix7642 : nand02 port map ( Y=>nx7643, A0=>nx4847, A1=>nx7859);
   ix7644 : inv01 port map ( Y=>nx7645, A=>nx4476);
   ix7646 : inv01 port map ( Y=>nx7647, A=>nx7645);
   ix7648 : inv01 port map ( Y=>nx7649, A=>nx4664);
   ix7650 : inv01 port map ( Y=>nx7651, A=>nx7649);
   ix7654 : nand02 port map ( Y=>nx7655, A0=>nx4894, A1=>nx7859);
   ix7656 : inv01 port map ( Y=>nx7657, A=>nx4860);
   ix7658 : inv01 port map ( Y=>nx7659, A=>nx7657);
   ix7660 : inv01 port map ( Y=>nx7661, A=>nx5048);
   ix7662 : inv01 port map ( Y=>nx7663, A=>nx7661);
   ix7666 : nand02 port map ( Y=>nx7667, A0=>nx4937, A1=>nx7859);
   ix7668 : inv01 port map ( Y=>nx7669, A=>nx5258);
   ix7670 : inv01 port map ( Y=>nx7671, A=>nx7669);
   ix7672 : inv01 port map ( Y=>nx7673, A=>nx5446);
   ix7674 : inv01 port map ( Y=>nx7675, A=>nx7673);
   ix7678 : nand02 port map ( Y=>nx7679, A0=>nx4985, A1=>nx7859);
   ix7680 : inv01 port map ( Y=>nx7681, A=>nx5642);
   ix7682 : inv01 port map ( Y=>nx7683, A=>nx7681);
   ix7684 : inv01 port map ( Y=>nx7685, A=>nx5830);
   ix7686 : inv01 port map ( Y=>nx7687, A=>nx7685);
   ix7690 : nand02 port map ( Y=>nx7691, A0=>nx5029, A1=>nx7859);
   ix7692 : inv01 port map ( Y=>nx7693, A=>nx6032);
   ix7694 : inv01 port map ( Y=>nx7695, A=>nx7693);
   ix7696 : inv01 port map ( Y=>nx7697, A=>nx6220);
   ix7698 : inv01 port map ( Y=>nx7699, A=>nx7697);
   ix7702 : nand02 port map ( Y=>nx7703, A0=>nx5075, A1=>nx7859);
   ix7704 : inv01 port map ( Y=>nx7705, A=>nx6416);
   ix7706 : inv01 port map ( Y=>nx7707, A=>nx7705);
   ix7708 : inv01 port map ( Y=>nx7709, A=>nx6604);
   ix7710 : inv01 port map ( Y=>nx7711, A=>nx7709);
   ix7714 : nand02 port map ( Y=>nx7715, A0=>nx5119, A1=>nx7861);
   ix7716 : inv01 port map ( Y=>nx7717, A=>nx6808);
   ix7718 : inv01 port map ( Y=>nx7719, A=>nx7717);
   ix7720 : inv01 port map ( Y=>nx7721, A=>nx6996);
   ix7722 : inv01 port map ( Y=>nx7723, A=>nx7721);
   ix7726 : nand02 port map ( Y=>nx7727, A0=>nx5165, A1=>nx7861);
   ix7728 : inv01 port map ( Y=>nx7729, A=>nx7192);
   ix7730 : inv01 port map ( Y=>nx7731, A=>nx7729);
   ix7732 : inv01 port map ( Y=>nx7733, A=>nx7380);
   ix7734 : inv01 port map ( Y=>nx7735, A=>nx7733);
   ix7736 : buf02 port map ( Y=>nx7737, A=>nx3523);
   ix7738 : buf02 port map ( Y=>nx7739, A=>nx3523);
   ix7740 : inv02 port map ( Y=>nx7741, A=>CNNIMGLOAD);
   ix7742 : inv02 port map ( Y=>nx7743, A=>CNNIMGLOAD);
   ix7744 : inv02 port map ( Y=>nx7745, A=>CNNIMGLOAD);
   ix7746 : inv02 port map ( Y=>nx7747, A=>CNNIMGLOAD);
   ix7748 : inv02 port map ( Y=>nx7749, A=>CNNIMGLOAD);
   ix7750 : inv02 port map ( Y=>nx7751, A=>CNNIMGLOAD);
   ix7752 : inv02 port map ( Y=>nx7753, A=>CNNIMGLOAD);
   ix7754 : inv02 port map ( Y=>nx7755, A=>CNNIMGLOAD);
   ix7756 : inv02 port map ( Y=>nx7757, A=>CNNIMGLOAD);
   ix7758 : inv02 port map ( Y=>nx7759, A=>CNNIMGLOAD);
   ix7760 : inv02 port map ( Y=>nx7761, A=>CNNIMGLOAD);
   ix7762 : inv02 port map ( Y=>nx7763, A=>CNNIMGLOAD);
   ix7764 : nor02_2x port map ( Y=>nx7765, A0=>nx3093, A1=>nx282);
   ix7766 : nor02_2x port map ( Y=>nx7767, A0=>nx3093, A1=>nx282);
   ix7768 : inv02 port map ( Y=>nx7769, A=>i8_reset1);
   ix7770 : inv02 port map ( Y=>nx7771, A=>i8_reset1);
   ix7772 : inv01 port map ( Y=>nx7773, A=>nx3921);
   ix7774 : inv02 port map ( Y=>nx7775, A=>nx7773);
   ix7776 : inv02 port map ( Y=>nx7777, A=>nx7773);
   ix7778 : inv02 port map ( Y=>nx7779, A=>nx7773);
   ix7780 : nor02_2x port map ( Y=>nx7781, A0=>nx3940, A1=>nx4126);
   ix7784 : inv02 port map ( Y=>nx7785, A=>nx7783);
   ix7786 : inv02 port map ( Y=>nx7787, A=>nx7783);
   ix7788 : inv02 port map ( Y=>nx7789, A=>nx7783);
   ix7790 : inv02 port map ( Y=>nx7791, A=>nx7783);
   ix7792 : inv02 port map ( Y=>nx7793, A=>nx7783);
   ix7794 : inv02 port map ( Y=>nx7795, A=>nx7783);
   ix7796 : inv02 port map ( Y=>nx7797, A=>nx7783);
   ix7798 : buf02 port map ( Y=>nx7799, A=>nx3971);
   ix7800 : buf02 port map ( Y=>nx7801, A=>nx3971);
   ix7802 : buf02 port map ( Y=>nx7803, A=>nx3999);
   ix7804 : buf02 port map ( Y=>nx7805, A=>nx3999);
   ix7806 : inv02 port map ( Y=>nx7807, A=>i8_counterout2_2);
   ix7808 : inv02 port map ( Y=>nx7809, A=>nx7913);
   ix7810 : nand02 port map ( Y=>nx7811, A0=>i8_reset2, A1=>zed);
   ix7812 : nor02_2x port map ( Y=>nx7813, A0=>i8_counterout2_0, A1=>
      i8_counterout2_1);
   ix7814 : inv02 port map ( Y=>nx7815, A=>i8_counterout2_3);
   ix7816 : inv02 port map ( Y=>nx7817, A=>i8_counterout2_3);
   ix7818 : inv02 port map ( Y=>nx7819, A=>i7_start);
   ix7820 : inv02 port map ( Y=>nx7821, A=>i7_start);
   ix7822 : inv02 port map ( Y=>nx7823, A=>i7_start);
   ix7824 : buf02 port map ( Y=>nx7825, A=>nx4246);
   ix7826 : buf02 port map ( Y=>nx7827, A=>nx4246);
   ix7828 : buf02 port map ( Y=>nx7829, A=>nx4271);
   ix7830 : buf02 port map ( Y=>nx7831, A=>nx4271);
   ix7832 : buf02 port map ( Y=>nx7833, A=>nx4274);
   ix7834 : buf02 port map ( Y=>nx7835, A=>nx4274);
   ix7836 : nor02_2x port map ( Y=>nx7837, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1);
   ix7838 : buf02 port map ( Y=>nx7839, A=>nx4303);
   ix7840 : buf02 port map ( Y=>nx7841, A=>nx4303);
   ix7842 : buf02 port map ( Y=>nx7843, A=>nx4405);
   ix7844 : buf02 port map ( Y=>nx7845, A=>nx4405);
   ix7846 : buf02 port map ( Y=>nx7847, A=>nx4407);
   ix7848 : buf02 port map ( Y=>nx7849, A=>nx4407);
   ix7852 : inv02 port map ( Y=>nx7853, A=>nx7851);
   ix7854 : inv02 port map ( Y=>nx7855, A=>nx7851);
   ix7856 : inv02 port map ( Y=>nx7857, A=>nx7851);
   ix7858 : inv02 port map ( Y=>nx7859, A=>nx7851);
   ix7860 : inv02 port map ( Y=>nx7861, A=>nx7851);
   ix7862 : nor02_2x port map ( Y=>nx7863, A0=>nx3940, A1=>i8_counterout2_1
   );
   ix7864 : nor02_2x port map ( Y=>nx7865, A0=>i8_counterout2_0, A1=>nx4126
   );
   ix7868 : inv02 port map ( Y=>nx7869, A=>nx7867);
   ix7870 : inv02 port map ( Y=>nx7871, A=>nx7867);
   ix7872 : inv02 port map ( Y=>nx7873, A=>nx7867);
   ix7874 : inv02 port map ( Y=>nx7875, A=>nx7867);
   ix7876 : inv02 port map ( Y=>nx7877, A=>i5_FAEN);
   ix7878 : inv02 port map ( Y=>nx7879, A=>i5_FAEN);
   ix7880 : inv02 port map ( Y=>nx7881, A=>i5_FAEN);
   ix7882 : inv02 port map ( Y=>nx7883, A=>i5_FAEN);
   ix7884 : inv02 port map ( Y=>nx7885, A=>i5_FAEN);
   ix7888 : inv02 port map ( Y=>nx7889, A=>nx7887);
   ix7890 : inv02 port map ( Y=>nx7891, A=>nx9398);
   ix7892 : inv02 port map ( Y=>nx7893, A=>nx9398);
   ix7894 : inv02 port map ( Y=>nx7895, A=>nx9398);
   ix7896 : inv02 port map ( Y=>nx7897, A=>nx9398);
   ix7898 : inv02 port map ( Y=>nx7899, A=>nx9398);
   ix7900 : inv02 port map ( Y=>nx7901, A=>nx9398);
   ix7906 : inv02 port map ( Y=>nx7907, A=>nx7959);
   ix7908 : inv02 port map ( Y=>nx7909, A=>nx7959);
   ix7910 : inv02 port map ( Y=>nx7911, A=>nx7807);
   ix7912 : inv02 port map ( Y=>nx7913, A=>nx7807);
   ix7956 : inv02 port map ( Y=>nx7957, A=>loadenable);
   ix7958 : inv02 port map ( Y=>nx7959, A=>loadenable);
   ix7960 : inv02 port map ( Y=>nx7961, A=>i8_counterout2_2);
   ix3524 : nor02_2x port map ( Y=>nx3523, A0=>nx66, A1=>Rst);
   ix69 : nor02_2x port map ( Y=>nx7399, A0=>nx8009, A1=>Rst);
   ix8008 : inv01 port map ( Y=>nx8009, A=>nx3565);
   ix3936 : nor02_2x port map ( Y=>nx3935, A0=>nx528, A1=>nx4151);
   ix3944 : nor02_2x port map ( Y=>nx3943, A0=>nx376, A1=>nx3940);
   ix3953 : nand02 port map ( Y=>nx7783, A0=>nx8011, A1=>nx7779);
   ix369 : aoi21 port map ( Y=>nx8011, A0=>i8_reset2, A1=>zed, B0=>nx4083);
   ix3158 : mux21 port map ( Y=>nx3157, A0=>nx8013, A1=>nx3967, S0=>nx7803);
   ix8012 : inv01 port map ( Y=>nx8013, A=>nx206);
   ix3178 : mux21 port map ( Y=>nx3177, A0=>nx8015, A1=>nx3979, S0=>nx7803);
   ix8014 : inv01 port map ( Y=>nx8015, A=>nx254);
   ix4014 : nor02_2x port map ( Y=>nx4013, A0=>nx3092, A1=>i8_counterout1_3
   );
   ix4030 : nor02_2x port map ( Y=>nx4029, A0=>nx314, A1=>nx7773);
   ix3148 : mux21 port map ( Y=>nx3147, A0=>nx8017, A1=>nx4033, S0=>nx7803);
   ix8016 : inv01 port map ( Y=>nx8017, A=>nx182);
   ix3168 : mux21 port map ( Y=>nx3167, A0=>nx8019, A1=>nx4050, S0=>nx7803);
   ix8018 : inv01 port map ( Y=>nx8019, A=>nx230);
   ix4067 : xnor2 port map ( Y=>nx4066, A0=>nx4059, A1=>nx8021);
   ix4070 : nand02 port map ( Y=>nx8021, A0=>nx8023, A1=>nx3979);
   ix8022 : inv01 port map ( Y=>nx8023, A=>nx3097);
   ix4080 : nor02_2x port map ( Y=>nx4079, A0=>nx3095, A1=>i8_counterout1_5
   );
   ix397 : xnor2 port map ( Y=>nx396, A0=>nx3940, A1=>nx4126);
   ix445 : xnor2 port map ( Y=>nx444, A0=>nx4151, A1=>nx8025);
   ix8024 : inv01 port map ( Y=>nx8025, A=>nx3101);
   ix481 : xnor2 port map ( Y=>nx480, A0=>nx4167, A1=>nx8027);
   ix8026 : inv01 port map ( Y=>nx8027, A=>nx458);
   ix465 : xnor2 port map ( Y=>nx464, A0=>nx4159, A1=>nx8029);
   ix8028 : inv01 port map ( Y=>nx8029, A=>nx3100);
   ix495 : xnor2 port map ( Y=>nx494, A0=>nx4177, A1=>nx8031);
   ix493 : nor02_2x port map ( Y=>nx8031, A0=>nx8033, A1=>i8_counterout2_6);
   ix4176 : nand02 port map ( Y=>nx8033, A0=>nx8029, A1=>nx4159);
   ix4199 : nor02_2x port map ( Y=>nx4198, A0=>nx602, A1=>nx7773);
   ix725 : xnor2 port map ( Y=>nx724, A0=>nx4283, A1=>nx8035);
   ix8034 : inv01 port map ( Y=>nx8035, A=>nx3111);
   ix4299 : nor02_2x port map ( Y=>nx4298, A0=>nx654, A1=>nx4309);
   ix4304 : nor02_2x port map ( Y=>nx4303, A0=>nx648, A1=>i7_start);
   ix675 : xnor2 port map ( Y=>nx674, A0=>nx4309, A1=>nx4317);
   ix709 : xnor2 port map ( Y=>nx708, A0=>nx4318, A1=>nx8037);
   ix703 : nor03_2x port map ( Y=>nx8037, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1, A2=>i7_counterout2_2);
   ix741 : xnor2 port map ( Y=>nx740, A0=>nx4333, A1=>nx8039);
   ix8038 : inv01 port map ( Y=>nx8039, A=>nx3109);
   ix759 : xnor2 port map ( Y=>nx758, A0=>nx4345, A1=>nx8041);
   ix8040 : inv01 port map ( Y=>nx8041, A=>nx3107);
   ix773 : xnor2 port map ( Y=>nx772, A0=>nx4355, A1=>nx8043);
   ix771 : nor02_2x port map ( Y=>nx8043, A0=>nx8045, A1=>i7_counterout2_6);
   ix4366 : nand02 port map ( Y=>nx8045, A0=>nx8039, A1=>nx4333);
   ix897 : nand03 port map ( Y=>nx4383, A0=>DataBus(12), A1=>DataBus(11), A2
      =>nx8047);
   ix8046 : inv01 port map ( Y=>nx8047, A=>nx4379);
   ix4387 : nor02_2x port map ( Y=>nx4386, A0=>nx3117, A1=>i7_counterout1_4
   );
   ix4408 : nor02_2x port map ( Y=>nx4407, A0=>nx856, A1=>i7_start);
   ix4420 : nor02_2x port map ( Y=>nx4419, A0=>nx3118, A1=>i7_counterout1_3
   );
   ix4438 : nor02_2x port map ( Y=>nx4437, A0=>nx3116, A1=>i7_counterout1_5
   );
   ix4463 : nor02_2x port map ( Y=>nx4462, A0=>nx3115, A1=>i7_counterout1_6
   );
   ix1101 : xnor2 port map ( Y=>nx1100, A0=>nx4487, A1=>nx8049);
   ix1099 : nor02_2x port map ( Y=>nx8049, A0=>nx8051, A1=>i7_counterout1_6
   );
   ix8050 : inv01 port map ( Y=>nx8051, A=>nx4437);
   ix691 : xnor2 port map ( Y=>nx690, A0=>nx4239, A1=>nx8053);
   ix685 : nor02_2x port map ( Y=>nx8053, A0=>i7_counterout2_0, A1=>
      i7_counterout2_1);
   ix551 : nand03 port map ( Y=>nx7433, A0=>nx4191, A1=>nx8055, A2=>
      EnableReadingFromCPU2);
   ix8054 : inv01 port map ( Y=>nx8055, A=>DataBus(15));
   ix4530 : nand03 port map ( Y=>nx7851, A0=>nx3925, A1=>CNNIMGLOAD, A2=>
      nx9396);
   ix1399 : nor02_2x port map ( Y=>nx1398, A0=>nx7511, A1=>nx8057);
   ix8056 : inv01 port map ( Y=>nx8057, A=>nx1188);
   ix1411 : nor02_2x port map ( Y=>nx1410, A0=>nx7511, A1=>nx8059);
   ix8058 : inv01 port map ( Y=>nx8059, A=>nx1202);
   ix1423 : nor02_2x port map ( Y=>nx1422, A0=>nx7511, A1=>nx8061);
   ix8060 : inv01 port map ( Y=>nx8061, A=>nx1216);
   ix1435 : nor02_2x port map ( Y=>nx1434, A0=>nx7511, A1=>nx8063);
   ix8062 : inv01 port map ( Y=>nx8063, A=>nx1230);
   ix1447 : nor02_2x port map ( Y=>nx1446, A0=>nx7511, A1=>nx8065);
   ix8064 : inv01 port map ( Y=>nx8065, A=>nx1244);
   ix1459 : nor02_2x port map ( Y=>nx1458, A0=>nx7511, A1=>nx8067);
   ix8066 : inv01 port map ( Y=>nx8067, A=>nx1258);
   ix1471 : nor02_2x port map ( Y=>nx1470, A0=>nx7511, A1=>nx8069);
   ix8068 : inv01 port map ( Y=>nx8069, A=>nx1272);
   ix1483 : nor02_2x port map ( Y=>nx1482, A0=>nx1388, A1=>nx8071);
   ix8070 : inv01 port map ( Y=>nx8071, A=>nx1286);
   ix1495 : nor02_2x port map ( Y=>nx1494, A0=>nx1388, A1=>nx8073);
   ix8072 : inv01 port map ( Y=>nx8073, A=>nx1300);
   ix1507 : nor02_2x port map ( Y=>nx1506, A0=>nx1388, A1=>nx8075);
   ix8074 : inv01 port map ( Y=>nx8075, A=>nx1314);
   ix1519 : nor02_2x port map ( Y=>nx1518, A0=>nx1388, A1=>nx8077);
   ix8076 : inv01 port map ( Y=>nx8077, A=>nx1328);
   ix1531 : nor02_2x port map ( Y=>nx1530, A0=>nx1388, A1=>nx8079);
   ix8078 : inv01 port map ( Y=>nx8079, A=>nx1342);
   ix1543 : nor02_2x port map ( Y=>nx1542, A0=>nx1388, A1=>nx8081);
   ix8080 : inv01 port map ( Y=>nx8081, A=>nx1356);
   ix1555 : nor02_2x port map ( Y=>nx1554, A0=>nx1388, A1=>nx8083);
   ix8082 : inv01 port map ( Y=>nx8083, A=>nx1370);
   ix5312 : nand03 port map ( Y=>nx7867, A0=>nx4227, A1=>nx7741, A2=>nx9396
   );
   ix4445 : nand03 port map ( Y=>nx7633, A0=>nx8085, A1=>nx4283, A2=>nx8087
   );
   ix8084 : inv01 port map ( Y=>nx8085, A=>nx7845);
   ix8086 : inv01 port map ( Y=>nx8087, A=>nx7841);
   ix1651 : mux21 port map ( Y=>Address(0), A0=>nx7039, A1=>nx7037, S0=>
      nx9398);
   ix1635 : xnor2 port map ( Y=>nx1634, A0=>nx7885, A1=>nx8089);
   ix8088 : inv01 port map ( Y=>nx8089, A=>nx7072);
   ix7056 : nor02_2x port map ( Y=>NOT_nx814, A0=>nx812, A1=>i7_tmp);
   ix7073 : mux21 port map ( Y=>nx7072, A0=>i5_MARo_0, A1=>OuterAddress(0), 
      S0=>nx9400);
   ix7076 : nor02_2x port map ( Y=>nx7887, A0=>nx7095, A1=>loadenable);
   ix1673 : mux21 port map ( Y=>Address(1), A0=>nx7081, A1=>nx7079, S0=>
      nx9400);
   ix1701 : mux21 port map ( Y=>Address(2), A0=>nx7100, A1=>nx7098, S0=>
      nx9400);
   ix7108 : mux21 port map ( Y=>nx7107, A0=>i5_MARo_1, A1=>OuterAddress(1), 
      S0=>nx9400);
   ix1729 : mux21 port map ( Y=>Address(3), A0=>nx7117, A1=>nx7115, S0=>
      nx9400);
   ix7127 : mux21 port map ( Y=>nx7126, A0=>i5_MARo_2, A1=>OuterAddress(2), 
      S0=>nx9400);
   ix7130 : mux21 port map ( Y=>nx7129, A0=>i5_MARo_3, A1=>OuterAddress(3), 
      S0=>nx9400);
   ix1757 : mux21 port map ( Y=>Address(4), A0=>nx7139, A1=>nx7137, S0=>
      nx9402);
   ix7149 : mux21 port map ( Y=>nx7148, A0=>i5_MARo_4, A1=>OuterAddress(4), 
      S0=>nx9402);
   ix1785 : mux21 port map ( Y=>Address(5), A0=>nx7159, A1=>nx7157, S0=>
      nx9402);
   ix7170 : mux21 port map ( Y=>nx7169, A0=>i5_MARo_5, A1=>OuterAddress(5), 
      S0=>nx9402);
   ix1813 : mux21 port map ( Y=>Address(6), A0=>nx7181, A1=>nx7178, S0=>
      nx9402);
   ix1841 : mux21 port map ( Y=>Address(7), A0=>nx7199, A1=>nx7197, S0=>
      nx9402);
   ix7210 : mux21 port map ( Y=>nx7209, A0=>i5_MARo_6, A1=>OuterAddress(6), 
      S0=>nx9402);
   ix7212 : mux21 port map ( Y=>nx7211, A0=>i5_MARo_7, A1=>OuterAddress(7), 
      S0=>nx9404);
   ix1869 : mux21 port map ( Y=>Address(8), A0=>nx7223, A1=>nx7221, S0=>
      nx9404);
   ix7234 : mux21 port map ( Y=>nx7233, A0=>i5_MARo_8, A1=>OuterAddress(8), 
      S0=>nx9404);
   ix1897 : mux21 port map ( Y=>Address(9), A0=>nx7243, A1=>nx7241, S0=>
      nx9404);
   ix7254 : mux21 port map ( Y=>nx7253, A0=>i5_MARo_9, A1=>OuterAddress(9), 
      S0=>nx9404);
   ix1925 : mux21 port map ( Y=>Address(10), A0=>nx7265, A1=>nx7262, S0=>
      nx9404);
   ix1953 : mux21 port map ( Y=>Address(11), A0=>nx7279, A1=>nx7277, S0=>
      nx9404);
   ix7288 : mux21 port map ( Y=>nx7287, A0=>i5_MARo_10, A1=>OuterAddress(10), 
      S0=>nx9406);
   ix7290 : mux21 port map ( Y=>nx7289, A0=>i5_MARo_11, A1=>OuterAddress(11), 
      S0=>nx9406);
   ix1981 : mux21 port map ( Y=>Address(12), A0=>nx7301, A1=>nx7298, S0=>
      nx9406);
   ix7311 : mux21 port map ( Y=>nx7310, A0=>i5_MARo_12, A1=>OuterAddress(12), 
      S0=>nx9406);
   ix2009 : mux21 port map ( Y=>Address(13), A0=>nx7321, A1=>nx7319, S0=>
      nx9406);
   ix7331 : mux21 port map ( Y=>nx7330, A0=>i5_MARo_13, A1=>OuterAddress(13), 
      S0=>nx9406);
   ix2037 : mux21 port map ( Y=>Address(14), A0=>nx7341, A1=>nx7339, S0=>
      nx9406);
   ix2065 : mux21 port map ( Y=>Address(15), A0=>nx7356, A1=>nx7354, S0=>
      nx9408);
   ix7366 : mux21 port map ( Y=>nx7365, A0=>i5_MARo_14, A1=>OuterAddress(14), 
      S0=>nx9408);
   ix7368 : mux21 port map ( Y=>nx7367, A0=>i5_MARo_15, A1=>OuterAddress(15), 
      S0=>nx9408);
   i8_lat_reset1_u1 : latchr port map ( QB=>nx5, D=>i8_nx74, CLK=>nx298, R=>
      DecompressedData1(255));
   i8_lat_reset1_u2 : inv01 port map ( Y=>i8_reset1, A=>nx5);
   i8_lat_tmp_u1 : latchs_ni port map ( QB=>nx8093, D=>
      DecompressedData1(255), CLK=>nx536, S=>nx540);
   i8_lat_tmp_u2 : inv02 port map ( Y=>zed, A=>nx8093);
   i8_lat_tmp_u3 : buf02 port map ( Y=>nx3955, A=>nx8093);
   i7_lat_tmp_u1 : latchs_ni port map ( QB=>nx8096, D=>
      DecompressedData1(255), CLK=>nx1140, S=>nx1148);
   i7_lat_tmp_u2 : inv02 port map ( Y=>i7_tmp, A=>nx8096);
   i7_lat_tmp_u3 : buf02 port map ( Y=>nx4277, A=>nx8096);
   i7_r28_lat_q_0_u1 : latchr port map ( QB=>nx8099, D=>nx9280, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(0), A=>nx8099);
   i7_r28_lat_q_0_u3 : buf02 port map ( Y=>nx5695, A=>nx8099);
   i8_r1_lat_q_0_u1 : latchr port map ( QB=>nx8102, D=>nx2122, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(0), A=>nx8102);
   i8_r1_lat_q_0_u3 : buf02 port map ( Y=>nx5697, A=>nx8102);
   i7_r28_lat_q_1_u1 : latchr port map ( QB=>nx8105, D=>nx9294, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(1), A=>nx8105);
   i7_r28_lat_q_1_u3 : buf02 port map ( Y=>nx5700, A=>nx8105);
   i8_r1_lat_q_1_u1 : latchr port map ( QB=>nx8108, D=>nx2148, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(1), A=>nx8108);
   i8_r1_lat_q_1_u3 : buf02 port map ( Y=>nx5703, A=>nx8108);
   i7_r28_lat_q_2_u1 : latchr port map ( QB=>nx8111, D=>nx9304, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(2), A=>nx8111);
   i7_r28_lat_q_2_u3 : buf02 port map ( Y=>nx5707, A=>nx8111);
   i8_r1_lat_q_2_u1 : latchr port map ( QB=>nx8114, D=>nx2174, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(2), A=>nx8114);
   i8_r1_lat_q_2_u3 : buf02 port map ( Y=>nx5709, A=>nx8114);
   i7_r28_lat_q_3_u1 : latchr port map ( QB=>nx8117, D=>nx9314, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(3), A=>nx8117);
   i7_r28_lat_q_3_u3 : buf02 port map ( Y=>nx5712, A=>nx8117);
   i8_r1_lat_q_3_u1 : latchr port map ( QB=>nx8120, D=>nx2200, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(3), A=>nx8120);
   i8_r1_lat_q_3_u3 : buf02 port map ( Y=>nx5715, A=>nx8120);
   i7_r28_lat_q_4_u1 : latchr port map ( QB=>nx8123, D=>nx9324, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(4), A=>nx8123);
   i7_r28_lat_q_4_u3 : buf02 port map ( Y=>nx5719, A=>nx8123);
   i8_r1_lat_q_4_u1 : latchr port map ( QB=>nx8126, D=>nx2226, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(4), A=>nx8126);
   i8_r1_lat_q_4_u3 : buf02 port map ( Y=>nx5721, A=>nx8126);
   i7_r28_lat_q_5_u1 : latchr port map ( QB=>nx8129, D=>nx9332, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(5), A=>nx8129);
   i7_r28_lat_q_5_u3 : buf02 port map ( Y=>nx5724, A=>nx8129);
   i8_r1_lat_q_5_u1 : latchr port map ( QB=>nx8132, D=>nx2252, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(5), A=>nx8132);
   i8_r1_lat_q_5_u3 : buf02 port map ( Y=>nx5727, A=>nx8132);
   i7_r28_lat_q_6_u1 : latchr port map ( QB=>nx8135, D=>nx9336, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(6), A=>nx8135);
   i7_r28_lat_q_6_u3 : buf02 port map ( Y=>nx5731, A=>nx8135);
   i8_r1_lat_q_6_u1 : latchr port map ( QB=>nx8138, D=>nx2278, CLK=>nx9288, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(6), A=>nx8138);
   i8_r1_lat_q_6_u3 : buf02 port map ( Y=>nx5733, A=>nx8138);
   i7_r28_lat_q_7_u1 : latchr port map ( QB=>nx8141, D=>nx9340, CLK=>nx2080, 
      R=>DecompressedData1(255));
   i7_r28_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(7), A=>nx8141);
   i7_r28_lat_q_7_u3 : buf02 port map ( Y=>nx5736, A=>nx8141);
   i8_r1_lat_q_7_u1 : latchr port map ( QB=>nx8144, D=>nx2304, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(7), A=>nx8144);
   i8_r1_lat_q_7_u3 : buf02 port map ( Y=>nx5739, A=>nx8144);
   i7_r27_lat_q_0_u1 : latchr port map ( QB=>nx8147, D=>nx9280, CLK=>nx2320, 
      R=>DecompressedData1(255));
   i7_r27_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(8), A=>nx8147);
   i7_r27_lat_q_0_u3 : buf02 port map ( Y=>nx5743, A=>nx8147);
   i8_r1_lat_q_8_u1 : latchr port map ( QB=>nx8150, D=>nx2334, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(8), A=>nx8150);
   i8_r1_lat_q_8_u3 : buf02 port map ( Y=>nx5745, A=>nx8150);
   i7_r27_lat_q_1_u1 : latchr port map ( QB=>nx8153, D=>nx9294, CLK=>nx2320, 
      R=>DecompressedData1(255));
   i7_r27_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(9), A=>nx8153);
   i7_r27_lat_q_1_u3 : buf02 port map ( Y=>nx5748, A=>nx8153);
   i8_r1_lat_q_9_u1 : latchr port map ( QB=>nx8156, D=>nx2358, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(9), A=>nx8156);
   i8_r1_lat_q_9_u3 : buf02 port map ( Y=>nx5751, A=>nx8156);
   i7_r27_lat_q_2_u1 : latchr port map ( QB=>nx8159, D=>nx9304, CLK=>nx2320, 
      R=>DecompressedData1(255));
   i7_r27_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(10), A=>nx8159
   );
   i7_r27_lat_q_2_u3 : buf02 port map ( Y=>nx5755, A=>nx8159);
   i8_r1_lat_q_10_u1 : latchr port map ( QB=>nx8162, D=>nx2382, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(10), A=>nx8162
   );
   i8_r1_lat_q_10_u3 : buf02 port map ( Y=>nx5757, A=>nx8162);
   i7_r27_lat_q_3_u1 : latchr port map ( QB=>nx8165, D=>nx9314, CLK=>nx2320, 
      R=>DecompressedData1(255));
   i7_r27_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(11), A=>nx8165
   );
   i7_r27_lat_q_3_u3 : buf02 port map ( Y=>nx5760, A=>nx8165);
   i8_r1_lat_q_11_u1 : latchr port map ( QB=>nx8168, D=>nx2406, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(11), A=>nx8168
   );
   i8_r1_lat_q_11_u3 : buf02 port map ( Y=>nx5763, A=>nx8168);
   i7_r27_lat_q_4_u1 : latchr port map ( QB=>nx8171, D=>nx9324, CLK=>nx2320, 
      R=>DecompressedData1(255));
   i7_r27_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(12), A=>nx8171
   );
   i7_r27_lat_q_4_u3 : buf02 port map ( Y=>nx5767, A=>nx8171);
   i8_r1_lat_q_12_u1 : latchr port map ( QB=>nx8174, D=>nx2430, CLK=>nx9290, 
      R=>DecompressedData1(255));
   i8_r1_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(12), A=>nx8174
   );
   i8_r1_lat_q_12_u3 : buf02 port map ( Y=>nx5769, A=>nx8174);
   i7_r26_lat_q_0_u1 : latchr port map ( QB=>nx8177, D=>nx9280, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(16), A=>nx8177
   );
   i7_r26_lat_q_0_u3 : buf02 port map ( Y=>nx5785, A=>nx8177);
   i8_r2_lat_q_0_u1 : latchr port map ( QB=>nx8180, D=>nx2524, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(16), A=>nx8180);
   i8_r2_lat_q_0_u3 : buf02 port map ( Y=>nx5787, A=>nx8180);
   i7_r26_lat_q_1_u1 : latchr port map ( QB=>nx8183, D=>nx9294, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(17), A=>nx8183
   );
   i7_r26_lat_q_1_u3 : buf02 port map ( Y=>nx5791, A=>nx8183);
   i8_r2_lat_q_1_u1 : latchr port map ( QB=>nx8186, D=>nx2548, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(17), A=>nx8186);
   i8_r2_lat_q_1_u3 : buf02 port map ( Y=>nx5793, A=>nx8186);
   i7_r26_lat_q_2_u1 : latchr port map ( QB=>nx8189, D=>nx9304, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(18), A=>nx8189
   );
   i7_r26_lat_q_2_u3 : buf02 port map ( Y=>nx5796, A=>nx8189);
   i8_r2_lat_q_2_u1 : latchr port map ( QB=>nx8192, D=>nx2572, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(18), A=>nx8192);
   i8_r2_lat_q_2_u3 : buf02 port map ( Y=>nx5799, A=>nx8192);
   i7_r26_lat_q_3_u1 : latchr port map ( QB=>nx8195, D=>nx9314, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(19), A=>nx8195
   );
   i7_r26_lat_q_3_u3 : buf02 port map ( Y=>nx5803, A=>nx8195);
   i8_r2_lat_q_3_u1 : latchr port map ( QB=>nx8198, D=>nx2596, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(19), A=>nx8198);
   i8_r2_lat_q_3_u3 : buf02 port map ( Y=>nx5805, A=>nx8198);
   i7_r26_lat_q_4_u1 : latchr port map ( QB=>nx8201, D=>nx9324, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(20), A=>nx8201
   );
   i7_r26_lat_q_4_u3 : buf02 port map ( Y=>nx5808, A=>nx8201);
   i8_r2_lat_q_4_u1 : latchr port map ( QB=>nx8204, D=>nx2620, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(20), A=>nx8204);
   i8_r2_lat_q_4_u3 : buf02 port map ( Y=>nx5811, A=>nx8204);
   i7_r26_lat_q_5_u1 : latchr port map ( QB=>nx8207, D=>nx9332, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(21), A=>nx8207
   );
   i7_r26_lat_q_5_u3 : buf02 port map ( Y=>nx5815, A=>nx8207);
   i8_r2_lat_q_5_u1 : latchr port map ( QB=>nx8210, D=>nx2644, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(21), A=>nx8210);
   i8_r2_lat_q_5_u3 : buf02 port map ( Y=>nx5817, A=>nx8210);
   i7_r26_lat_q_6_u1 : latchr port map ( QB=>nx8213, D=>nx9336, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(22), A=>nx8213
   );
   i7_r26_lat_q_6_u3 : buf02 port map ( Y=>nx5820, A=>nx8213);
   i8_r2_lat_q_6_u1 : latchr port map ( QB=>nx8216, D=>nx2668, CLK=>nx9344, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(22), A=>nx8216);
   i8_r2_lat_q_6_u3 : buf02 port map ( Y=>nx5823, A=>nx8216);
   i7_r26_lat_q_7_u1 : latchr port map ( QB=>nx8219, D=>nx9340, CLK=>nx2494, 
      R=>DecompressedData1(255));
   i7_r26_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(23), A=>nx8219
   );
   i7_r26_lat_q_7_u3 : buf02 port map ( Y=>nx5827, A=>nx8219);
   i8_r2_lat_q_7_u1 : latchr port map ( QB=>nx8222, D=>nx2692, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(23), A=>nx8222);
   i8_r2_lat_q_7_u3 : buf02 port map ( Y=>nx5829, A=>nx8222);
   i7_r25_lat_q_0_u1 : latchr port map ( QB=>nx8225, D=>nx9280, CLK=>nx2708, 
      R=>DecompressedData1(255));
   i7_r25_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(24), A=>nx8225
   );
   i7_r25_lat_q_0_u3 : buf02 port map ( Y=>nx5833, A=>nx8225);
   i8_r2_lat_q_8_u1 : latchr port map ( QB=>nx8228, D=>nx2722, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(24), A=>nx8228);
   i8_r2_lat_q_8_u3 : buf02 port map ( Y=>nx5835, A=>nx8228);
   i7_r25_lat_q_1_u1 : latchr port map ( QB=>nx8231, D=>nx9294, CLK=>nx2708, 
      R=>DecompressedData1(255));
   i7_r25_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(25), A=>nx8231
   );
   i7_r25_lat_q_1_u3 : buf02 port map ( Y=>nx5838, A=>nx8231);
   i8_r2_lat_q_9_u1 : latchr port map ( QB=>nx8234, D=>nx2746, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(25), A=>nx8234);
   i8_r2_lat_q_9_u3 : buf02 port map ( Y=>nx5841, A=>nx8234);
   i7_r25_lat_q_2_u1 : latchr port map ( QB=>nx8237, D=>nx9304, CLK=>nx2708, 
      R=>DecompressedData1(255));
   i7_r25_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(26), A=>nx8237
   );
   i7_r25_lat_q_2_u3 : buf02 port map ( Y=>nx5845, A=>nx8237);
   i8_r2_lat_q_10_u1 : latchr port map ( QB=>nx8240, D=>nx2770, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(26), A=>nx8240
   );
   i8_r2_lat_q_10_u3 : buf02 port map ( Y=>nx5847, A=>nx8240);
   i7_r25_lat_q_3_u1 : latchr port map ( QB=>nx8243, D=>nx9314, CLK=>nx2708, 
      R=>DecompressedData1(255));
   i7_r25_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(27), A=>nx8243
   );
   i7_r25_lat_q_3_u3 : buf02 port map ( Y=>nx5850, A=>nx8243);
   i8_r2_lat_q_11_u1 : latchr port map ( QB=>nx8246, D=>nx2794, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(27), A=>nx8246
   );
   i8_r2_lat_q_11_u3 : buf02 port map ( Y=>nx5853, A=>nx8246);
   i7_r25_lat_q_4_u1 : latchr port map ( QB=>nx8249, D=>nx9324, CLK=>nx2708, 
      R=>DecompressedData1(255));
   i7_r25_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(28), A=>nx8249
   );
   i7_r25_lat_q_4_u3 : buf02 port map ( Y=>nx5857, A=>nx8249);
   i8_r2_lat_q_12_u1 : latchr port map ( QB=>nx8252, D=>nx2818, CLK=>nx9346, 
      R=>DecompressedData1(255));
   i8_r2_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(28), A=>nx8252
   );
   i8_r2_lat_q_12_u3 : buf02 port map ( Y=>nx5859, A=>nx8252);
   i7_r24_lat_q_0_u1 : latchr port map ( QB=>nx8255, D=>nx9280, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(32), A=>nx8255
   );
   i7_r24_lat_q_0_u3 : buf02 port map ( Y=>nx5875, A=>nx8255);
   i8_r3_lat_q_0_u1 : latchr port map ( QB=>nx8258, D=>nx2914, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(32), A=>nx8258);
   i8_r3_lat_q_0_u3 : buf02 port map ( Y=>nx5877, A=>nx8258);
   i7_r24_lat_q_1_u1 : latchr port map ( QB=>nx8261, D=>nx9294, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(33), A=>nx8261
   );
   i7_r24_lat_q_1_u3 : buf02 port map ( Y=>nx5881, A=>nx8261);
   i8_r3_lat_q_1_u1 : latchr port map ( QB=>nx8264, D=>nx2938, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(33), A=>nx8264);
   i8_r3_lat_q_1_u3 : buf02 port map ( Y=>nx5883, A=>nx8264);
   i7_r24_lat_q_2_u1 : latchr port map ( QB=>nx8267, D=>nx9304, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(34), A=>nx8267
   );
   i7_r24_lat_q_2_u3 : buf02 port map ( Y=>nx5886, A=>nx8267);
   i8_r3_lat_q_2_u1 : latchr port map ( QB=>nx8270, D=>nx2962, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(34), A=>nx8270);
   i8_r3_lat_q_2_u3 : buf02 port map ( Y=>nx5889, A=>nx8270);
   i7_r24_lat_q_3_u1 : latchr port map ( QB=>nx8273, D=>nx9314, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(35), A=>nx8273
   );
   i7_r24_lat_q_3_u3 : buf02 port map ( Y=>nx5893, A=>nx8273);
   i8_r3_lat_q_3_u1 : latchr port map ( QB=>nx8276, D=>nx2986, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(35), A=>nx8276);
   i8_r3_lat_q_3_u3 : buf02 port map ( Y=>nx5895, A=>nx8276);
   i7_r24_lat_q_4_u1 : latchr port map ( QB=>nx8279, D=>nx9324, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(36), A=>nx8279
   );
   i7_r24_lat_q_4_u3 : buf02 port map ( Y=>nx5898, A=>nx8279);
   i8_r3_lat_q_4_u1 : latchr port map ( QB=>nx8282, D=>nx3010, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(36), A=>nx8282);
   i8_r3_lat_q_4_u3 : buf02 port map ( Y=>nx5901, A=>nx8282);
   i7_r24_lat_q_5_u1 : latchr port map ( QB=>nx8285, D=>nx9332, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(37), A=>nx8285
   );
   i7_r24_lat_q_5_u3 : buf02 port map ( Y=>nx5905, A=>nx8285);
   i8_r3_lat_q_5_u1 : latchr port map ( QB=>nx8288, D=>nx3034, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(37), A=>nx8288);
   i8_r3_lat_q_5_u3 : buf02 port map ( Y=>nx5907, A=>nx8288);
   i7_r24_lat_q_6_u1 : latchr port map ( QB=>nx8291, D=>nx9336, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(38), A=>nx8291
   );
   i7_r24_lat_q_6_u3 : buf02 port map ( Y=>nx5910, A=>nx8291);
   i8_r3_lat_q_6_u1 : latchr port map ( QB=>nx8294, D=>nx3058, CLK=>nx9348, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(38), A=>nx8294);
   i8_r3_lat_q_6_u3 : buf02 port map ( Y=>nx5913, A=>nx8294);
   i7_r24_lat_q_7_u1 : latchr port map ( QB=>nx8297, D=>nx9340, CLK=>nx2888, 
      R=>DecompressedData1(255));
   i7_r24_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(39), A=>nx8297
   );
   i7_r24_lat_q_7_u3 : buf02 port map ( Y=>nx5917, A=>nx8297);
   i8_r3_lat_q_7_u1 : latchr port map ( QB=>nx8300, D=>nx3082, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(39), A=>nx8300);
   i8_r3_lat_q_7_u3 : buf02 port map ( Y=>nx5919, A=>nx8300);
   i7_r23_lat_q_0_u1 : latchr port map ( QB=>nx8303, D=>nx9280, CLK=>nx3098, 
      R=>DecompressedData1(255));
   i7_r23_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(40), A=>nx8303
   );
   i7_r23_lat_q_0_u3 : buf02 port map ( Y=>nx5922, A=>nx8303);
   i8_r3_lat_q_8_u1 : latchr port map ( QB=>nx8306, D=>nx3112, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(40), A=>nx8306);
   i8_r3_lat_q_8_u3 : buf02 port map ( Y=>nx5925, A=>nx8306);
   i7_r23_lat_q_1_u1 : latchr port map ( QB=>nx8309, D=>nx9294, CLK=>nx3098, 
      R=>DecompressedData1(255));
   i7_r23_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(41), A=>nx8309
   );
   i7_r23_lat_q_1_u3 : buf02 port map ( Y=>nx5929, A=>nx8309);
   i8_r3_lat_q_9_u1 : latchr port map ( QB=>nx8312, D=>nx3136, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(41), A=>nx8312);
   i8_r3_lat_q_9_u3 : buf02 port map ( Y=>nx5931, A=>nx8312);
   i7_r23_lat_q_2_u1 : latchr port map ( QB=>nx8315, D=>nx9304, CLK=>nx3098, 
      R=>DecompressedData1(255));
   i7_r23_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(42), A=>nx8315
   );
   i7_r23_lat_q_2_u3 : buf02 port map ( Y=>nx5934, A=>nx8315);
   i8_r3_lat_q_10_u1 : latchr port map ( QB=>nx8318, D=>nx3160, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(42), A=>nx8318
   );
   i8_r3_lat_q_10_u3 : buf02 port map ( Y=>nx5937, A=>nx8318);
   i7_r23_lat_q_3_u1 : latchr port map ( QB=>nx8321, D=>nx9314, CLK=>nx3098, 
      R=>DecompressedData1(255));
   i7_r23_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(43), A=>nx8321
   );
   i7_r23_lat_q_3_u3 : buf02 port map ( Y=>nx5941, A=>nx8321);
   i8_r3_lat_q_11_u1 : latchr port map ( QB=>nx8324, D=>nx3184, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(43), A=>nx8324
   );
   i8_r3_lat_q_11_u3 : buf02 port map ( Y=>nx5943, A=>nx8324);
   i7_r23_lat_q_4_u1 : latchr port map ( QB=>nx8327, D=>nx9324, CLK=>nx3098, 
      R=>DecompressedData1(255));
   i7_r23_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(44), A=>nx8327
   );
   i7_r23_lat_q_4_u3 : buf02 port map ( Y=>nx5946, A=>nx8327);
   i8_r3_lat_q_12_u1 : latchr port map ( QB=>nx8330, D=>nx3208, CLK=>nx9350, 
      R=>DecompressedData1(255));
   i8_r3_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(44), A=>nx8330
   );
   i8_r3_lat_q_12_u3 : buf02 port map ( Y=>nx5949, A=>nx8330);
   i7_r22_lat_q_0_u1 : latchr port map ( QB=>nx8333, D=>nx9280, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(48), A=>nx8333
   );
   i7_r22_lat_q_0_u3 : buf02 port map ( Y=>nx5965, A=>nx8333);
   i8_r4_lat_q_0_u1 : latchr port map ( QB=>nx8336, D=>nx3302, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(48), A=>nx8336);
   i8_r4_lat_q_0_u3 : buf02 port map ( Y=>nx5967, A=>nx8336);
   i7_r22_lat_q_1_u1 : latchr port map ( QB=>nx8339, D=>nx9294, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(49), A=>nx8339
   );
   i7_r22_lat_q_1_u3 : buf02 port map ( Y=>nx5970, A=>nx8339);
   i8_r4_lat_q_1_u1 : latchr port map ( QB=>nx8342, D=>nx3326, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(49), A=>nx8342);
   i8_r4_lat_q_1_u3 : buf02 port map ( Y=>nx5973, A=>nx8342);
   i7_r22_lat_q_2_u1 : latchr port map ( QB=>nx8345, D=>nx9304, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(50), A=>nx8345
   );
   i7_r22_lat_q_2_u3 : buf02 port map ( Y=>nx5977, A=>nx8345);
   i8_r4_lat_q_2_u1 : latchr port map ( QB=>nx8348, D=>nx3350, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(50), A=>nx8348);
   i8_r4_lat_q_2_u3 : buf02 port map ( Y=>nx5979, A=>nx8348);
   i7_r22_lat_q_3_u1 : latchr port map ( QB=>nx8351, D=>nx9314, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(51), A=>nx8351
   );
   i7_r22_lat_q_3_u3 : buf02 port map ( Y=>nx5982, A=>nx8351);
   i8_r4_lat_q_3_u1 : latchr port map ( QB=>nx8354, D=>nx3374, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(51), A=>nx8354);
   i8_r4_lat_q_3_u3 : buf02 port map ( Y=>nx5985, A=>nx8354);
   i7_r22_lat_q_4_u1 : latchr port map ( QB=>nx8357, D=>nx9324, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(52), A=>nx8357
   );
   i7_r22_lat_q_4_u3 : buf02 port map ( Y=>nx5989, A=>nx8357);
   i8_r4_lat_q_4_u1 : latchr port map ( QB=>nx8360, D=>nx3398, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(52), A=>nx8360);
   i8_r4_lat_q_4_u3 : buf02 port map ( Y=>nx5991, A=>nx8360);
   i7_r22_lat_q_5_u1 : latchr port map ( QB=>nx8363, D=>nx9332, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(53), A=>nx8363
   );
   i7_r22_lat_q_5_u3 : buf02 port map ( Y=>nx5994, A=>nx8363);
   i8_r4_lat_q_5_u1 : latchr port map ( QB=>nx8366, D=>nx3422, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(53), A=>nx8366);
   i8_r4_lat_q_5_u3 : buf02 port map ( Y=>nx5997, A=>nx8366);
   i7_r22_lat_q_6_u1 : latchr port map ( QB=>nx8369, D=>nx9336, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(54), A=>nx8369
   );
   i7_r22_lat_q_6_u3 : buf02 port map ( Y=>nx6001, A=>nx8369);
   i8_r4_lat_q_6_u1 : latchr port map ( QB=>nx8372, D=>nx3446, CLK=>nx9352, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(54), A=>nx8372);
   i8_r4_lat_q_6_u3 : buf02 port map ( Y=>nx6003, A=>nx8372);
   i7_r22_lat_q_7_u1 : latchr port map ( QB=>nx8375, D=>nx9340, CLK=>nx3272, 
      R=>DecompressedData1(255));
   i7_r22_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(55), A=>nx8375
   );
   i7_r22_lat_q_7_u3 : buf02 port map ( Y=>nx6007, A=>nx8375);
   i8_r4_lat_q_7_u1 : latchr port map ( QB=>nx8378, D=>nx3470, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(55), A=>nx8378);
   i8_r4_lat_q_7_u3 : buf02 port map ( Y=>nx6009, A=>nx8378);
   i7_r21_lat_q_0_u1 : latchr port map ( QB=>nx8381, D=>nx9282, CLK=>nx3486, 
      R=>DecompressedData1(255));
   i7_r21_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(56), A=>nx8381
   );
   i7_r21_lat_q_0_u3 : buf02 port map ( Y=>nx6013, A=>nx8381);
   i8_r4_lat_q_8_u1 : latchr port map ( QB=>nx8384, D=>nx3500, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(56), A=>nx8384);
   i8_r4_lat_q_8_u3 : buf02 port map ( Y=>nx6015, A=>nx8384);
   i7_r21_lat_q_1_u1 : latchr port map ( QB=>nx8387, D=>nx9296, CLK=>nx3486, 
      R=>DecompressedData1(255));
   i7_r21_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(57), A=>nx8387
   );
   i7_r21_lat_q_1_u3 : buf02 port map ( Y=>nx6018, A=>nx8387);
   i8_r4_lat_q_9_u1 : latchr port map ( QB=>nx8390, D=>nx3524, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(57), A=>nx8390);
   i8_r4_lat_q_9_u3 : buf02 port map ( Y=>nx6021, A=>nx8390);
   i7_r21_lat_q_2_u1 : latchr port map ( QB=>nx8393, D=>nx9306, CLK=>nx3486, 
      R=>DecompressedData1(255));
   i7_r21_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(58), A=>nx8393
   );
   i7_r21_lat_q_2_u3 : buf02 port map ( Y=>nx6025, A=>nx8393);
   i8_r4_lat_q_10_u1 : latchr port map ( QB=>nx8396, D=>nx3548, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(58), A=>nx8396
   );
   i8_r4_lat_q_10_u3 : buf02 port map ( Y=>nx6027, A=>nx8396);
   i7_r21_lat_q_3_u1 : latchr port map ( QB=>nx8399, D=>nx9316, CLK=>nx3486, 
      R=>DecompressedData1(255));
   i7_r21_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(59), A=>nx8399
   );
   i7_r21_lat_q_3_u3 : buf02 port map ( Y=>nx6031, A=>nx8399);
   i8_r4_lat_q_11_u1 : latchr port map ( QB=>nx8402, D=>nx3572, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(59), A=>nx8402
   );
   i8_r4_lat_q_11_u3 : buf02 port map ( Y=>nx6033, A=>nx8402);
   i7_r21_lat_q_4_u1 : latchr port map ( QB=>nx8405, D=>nx9326, CLK=>nx3486, 
      R=>DecompressedData1(255));
   i7_r21_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(60), A=>nx8405
   );
   i7_r21_lat_q_4_u3 : buf02 port map ( Y=>nx6037, A=>nx8405);
   i8_r4_lat_q_12_u1 : latchr port map ( QB=>nx8408, D=>nx3596, CLK=>nx9354, 
      R=>DecompressedData1(255));
   i8_r4_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(60), A=>nx8408
   );
   i8_r4_lat_q_12_u3 : buf02 port map ( Y=>nx6039, A=>nx8408);
   i7_r20_lat_q_0_u1 : latchr port map ( QB=>nx8411, D=>nx9282, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(64), A=>nx8411
   );
   i7_r20_lat_q_0_u3 : buf02 port map ( Y=>nx6055, A=>nx8411);
   i8_r5_lat_q_0_u1 : latchr port map ( QB=>nx8414, D=>nx3702, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(64), A=>nx8414);
   i8_r5_lat_q_0_u3 : buf02 port map ( Y=>nx6057, A=>nx8414);
   i7_r20_lat_q_1_u1 : latchr port map ( QB=>nx8417, D=>nx9296, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(65), A=>nx8417
   );
   i7_r20_lat_q_1_u3 : buf02 port map ( Y=>nx6061, A=>nx8417);
   i8_r5_lat_q_1_u1 : latchr port map ( QB=>nx8420, D=>nx3726, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(65), A=>nx8420);
   i8_r5_lat_q_1_u3 : buf02 port map ( Y=>nx6063, A=>nx8420);
   i7_r20_lat_q_2_u1 : latchr port map ( QB=>nx8423, D=>nx9306, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(66), A=>nx8423
   );
   i7_r20_lat_q_2_u3 : buf02 port map ( Y=>nx6066, A=>nx8423);
   i8_r5_lat_q_2_u1 : latchr port map ( QB=>nx8426, D=>nx3750, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(66), A=>nx8426);
   i8_r5_lat_q_2_u3 : buf02 port map ( Y=>nx6069, A=>nx8426);
   i7_r20_lat_q_3_u1 : latchr port map ( QB=>nx8429, D=>nx9316, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(67), A=>nx8429
   );
   i7_r20_lat_q_3_u3 : buf02 port map ( Y=>nx6073, A=>nx8429);
   i8_r5_lat_q_3_u1 : latchr port map ( QB=>nx8432, D=>nx3774, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(67), A=>nx8432);
   i8_r5_lat_q_3_u3 : buf02 port map ( Y=>nx6075, A=>nx8432);
   i7_r20_lat_q_4_u1 : latchr port map ( QB=>nx8435, D=>nx9326, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(68), A=>nx8435
   );
   i7_r20_lat_q_4_u3 : buf02 port map ( Y=>nx6078, A=>nx8435);
   i8_r5_lat_q_4_u1 : latchr port map ( QB=>nx8438, D=>nx3798, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(68), A=>nx8438);
   i8_r5_lat_q_4_u3 : buf02 port map ( Y=>nx6081, A=>nx8438);
   i7_r20_lat_q_5_u1 : latchr port map ( QB=>nx8441, D=>nx9332, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(69), A=>nx8441
   );
   i7_r20_lat_q_5_u3 : buf02 port map ( Y=>nx6085, A=>nx8441);
   i8_r5_lat_q_5_u1 : latchr port map ( QB=>nx8444, D=>nx3822, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(69), A=>nx8444);
   i8_r5_lat_q_5_u3 : buf02 port map ( Y=>nx6087, A=>nx8444);
   i7_r20_lat_q_6_u1 : latchr port map ( QB=>nx8447, D=>nx9336, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(70), A=>nx8447
   );
   i7_r20_lat_q_6_u3 : buf02 port map ( Y=>nx6090, A=>nx8447);
   i8_r5_lat_q_6_u1 : latchr port map ( QB=>nx8450, D=>nx3846, CLK=>nx9356, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(70), A=>nx8450);
   i8_r5_lat_q_6_u3 : buf02 port map ( Y=>nx6093, A=>nx8450);
   i7_r20_lat_q_7_u1 : latchr port map ( QB=>nx8453, D=>nx9340, CLK=>nx3668, 
      R=>DecompressedData1(255));
   i7_r20_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(71), A=>nx8453
   );
   i7_r20_lat_q_7_u3 : buf02 port map ( Y=>nx6097, A=>nx8453);
   i8_r5_lat_q_7_u1 : latchr port map ( QB=>nx8456, D=>nx3870, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(71), A=>nx8456);
   i8_r5_lat_q_7_u3 : buf02 port map ( Y=>nx6099, A=>nx8456);
   i7_r19_lat_q_0_u1 : latchr port map ( QB=>nx8459, D=>nx9282, CLK=>nx3886, 
      R=>DecompressedData1(255));
   i7_r19_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(72), A=>nx8459
   );
   i7_r19_lat_q_0_u3 : buf02 port map ( Y=>nx6102, A=>nx8459);
   i8_r5_lat_q_8_u1 : latchr port map ( QB=>nx8462, D=>nx3900, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(72), A=>nx8462);
   i8_r5_lat_q_8_u3 : buf02 port map ( Y=>nx6105, A=>nx8462);
   i7_r19_lat_q_1_u1 : latchr port map ( QB=>nx8465, D=>nx9296, CLK=>nx3886, 
      R=>DecompressedData1(255));
   i7_r19_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(73), A=>nx8465
   );
   i7_r19_lat_q_1_u3 : buf02 port map ( Y=>nx6109, A=>nx8465);
   i8_r5_lat_q_9_u1 : latchr port map ( QB=>nx8468, D=>nx3924, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(73), A=>nx8468);
   i8_r5_lat_q_9_u3 : buf02 port map ( Y=>nx6111, A=>nx8468);
   i7_r19_lat_q_2_u1 : latchr port map ( QB=>nx8471, D=>nx9306, CLK=>nx3886, 
      R=>DecompressedData1(255));
   i7_r19_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(74), A=>nx8471
   );
   i7_r19_lat_q_2_u3 : buf02 port map ( Y=>nx6114, A=>nx8471);
   i8_r5_lat_q_10_u1 : latchr port map ( QB=>nx8474, D=>nx3948, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(74), A=>nx8474
   );
   i8_r5_lat_q_10_u3 : buf02 port map ( Y=>nx6117, A=>nx8474);
   i7_r19_lat_q_3_u1 : latchr port map ( QB=>nx8477, D=>nx9316, CLK=>nx3886, 
      R=>DecompressedData1(255));
   i7_r19_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(75), A=>nx8477
   );
   i7_r19_lat_q_3_u3 : buf02 port map ( Y=>nx6121, A=>nx8477);
   i8_r5_lat_q_11_u1 : latchr port map ( QB=>nx8480, D=>nx3972, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(75), A=>nx8480
   );
   i8_r5_lat_q_11_u3 : buf02 port map ( Y=>nx6123, A=>nx8480);
   i7_r19_lat_q_4_u1 : latchr port map ( QB=>nx8483, D=>nx9326, CLK=>nx3886, 
      R=>DecompressedData1(255));
   i7_r19_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(76), A=>nx8483
   );
   i7_r19_lat_q_4_u3 : buf02 port map ( Y=>nx6126, A=>nx8483);
   i8_r5_lat_q_12_u1 : latchr port map ( QB=>nx8486, D=>nx3996, CLK=>nx9358, 
      R=>DecompressedData1(255));
   i8_r5_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(76), A=>nx8486
   );
   i8_r5_lat_q_12_u3 : buf02 port map ( Y=>nx6129, A=>nx8486);
   i7_r18_lat_q_0_u1 : latchr port map ( QB=>nx8489, D=>nx9282, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(80), A=>nx8489
   );
   i7_r18_lat_q_0_u3 : buf02 port map ( Y=>nx6145, A=>nx8489);
   i8_r6_lat_q_0_u1 : latchr port map ( QB=>nx8492, D=>nx4086, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(80), A=>nx8492);
   i8_r6_lat_q_0_u3 : buf02 port map ( Y=>nx6147, A=>nx8492);
   i7_r18_lat_q_1_u1 : latchr port map ( QB=>nx8495, D=>nx9296, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(81), A=>nx8495
   );
   i7_r18_lat_q_1_u3 : buf02 port map ( Y=>nx6150, A=>nx8495);
   i8_r6_lat_q_1_u1 : latchr port map ( QB=>nx8498, D=>nx4110, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(81), A=>nx8498);
   i8_r6_lat_q_1_u3 : buf02 port map ( Y=>nx6153, A=>nx8498);
   i7_r18_lat_q_2_u1 : latchr port map ( QB=>nx8501, D=>nx9306, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(82), A=>nx8501
   );
   i7_r18_lat_q_2_u3 : buf02 port map ( Y=>nx6157, A=>nx8501);
   i8_r6_lat_q_2_u1 : latchr port map ( QB=>nx8504, D=>nx4134, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(82), A=>nx8504);
   i8_r6_lat_q_2_u3 : buf02 port map ( Y=>nx6159, A=>nx8504);
   i7_r18_lat_q_3_u1 : latchr port map ( QB=>nx8507, D=>nx9316, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(83), A=>nx8507
   );
   i7_r18_lat_q_3_u3 : buf02 port map ( Y=>nx6162, A=>nx8507);
   i8_r6_lat_q_3_u1 : latchr port map ( QB=>nx8510, D=>nx4158, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(83), A=>nx8510);
   i8_r6_lat_q_3_u3 : buf02 port map ( Y=>nx6165, A=>nx8510);
   i7_r18_lat_q_4_u1 : latchr port map ( QB=>nx8513, D=>nx9326, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(84), A=>nx8513
   );
   i7_r18_lat_q_4_u3 : buf02 port map ( Y=>nx6169, A=>nx8513);
   i8_r6_lat_q_4_u1 : latchr port map ( QB=>nx8516, D=>nx4182, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(84), A=>nx8516);
   i8_r6_lat_q_4_u3 : buf02 port map ( Y=>nx6171, A=>nx8516);
   i7_r18_lat_q_5_u1 : latchr port map ( QB=>nx8519, D=>nx9332, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(85), A=>nx8519
   );
   i7_r18_lat_q_5_u3 : buf02 port map ( Y=>nx6174, A=>nx8519);
   i8_r6_lat_q_5_u1 : latchr port map ( QB=>nx8522, D=>nx4206, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(85), A=>nx8522);
   i8_r6_lat_q_5_u3 : buf02 port map ( Y=>nx6177, A=>nx8522);
   i7_r18_lat_q_6_u1 : latchr port map ( QB=>nx8525, D=>nx9336, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(86), A=>nx8525
   );
   i7_r18_lat_q_6_u3 : buf02 port map ( Y=>nx6181, A=>nx8525);
   i8_r6_lat_q_6_u1 : latchr port map ( QB=>nx8528, D=>nx4230, CLK=>nx9360, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(86), A=>nx8528);
   i8_r6_lat_q_6_u3 : buf02 port map ( Y=>nx6183, A=>nx8528);
   i7_r18_lat_q_7_u1 : latchr port map ( QB=>nx8531, D=>nx9340, CLK=>nx4060, 
      R=>DecompressedData1(255));
   i7_r18_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(87), A=>nx8531
   );
   i7_r18_lat_q_7_u3 : buf02 port map ( Y=>nx6186, A=>nx8531);
   i8_r6_lat_q_7_u1 : latchr port map ( QB=>nx8534, D=>nx4254, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(87), A=>nx8534);
   i8_r6_lat_q_7_u3 : buf02 port map ( Y=>nx6189, A=>nx8534);
   i7_r17_lat_q_0_u1 : latchr port map ( QB=>nx8537, D=>nx9282, CLK=>nx4270, 
      R=>DecompressedData1(255));
   i7_r17_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(88), A=>nx8537
   );
   i7_r17_lat_q_0_u3 : buf02 port map ( Y=>nx6193, A=>nx8537);
   i8_r6_lat_q_8_u1 : latchr port map ( QB=>nx8540, D=>nx4284, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(88), A=>nx8540);
   i8_r6_lat_q_8_u3 : buf02 port map ( Y=>nx6195, A=>nx8540);
   i7_r17_lat_q_1_u1 : latchr port map ( QB=>nx8543, D=>nx9296, CLK=>nx4270, 
      R=>DecompressedData1(255));
   i7_r17_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(89), A=>nx8543
   );
   i7_r17_lat_q_1_u3 : buf02 port map ( Y=>nx6198, A=>nx8543);
   i8_r6_lat_q_9_u1 : latchr port map ( QB=>nx8546, D=>nx4308, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(89), A=>nx8546);
   i8_r6_lat_q_9_u3 : buf02 port map ( Y=>nx6201, A=>nx8546);
   i7_r17_lat_q_2_u1 : latchr port map ( QB=>nx8549, D=>nx9306, CLK=>nx4270, 
      R=>DecompressedData1(255));
   i7_r17_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(90), A=>nx8549
   );
   i7_r17_lat_q_2_u3 : buf02 port map ( Y=>nx6205, A=>nx8549);
   i8_r6_lat_q_10_u1 : latchr port map ( QB=>nx8552, D=>nx4332, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(90), A=>nx8552
   );
   i8_r6_lat_q_10_u3 : buf02 port map ( Y=>nx6207, A=>nx8552);
   i7_r17_lat_q_3_u1 : latchr port map ( QB=>nx8555, D=>nx9316, CLK=>nx4270, 
      R=>DecompressedData1(255));
   i7_r17_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(91), A=>nx8555
   );
   i7_r17_lat_q_3_u3 : buf02 port map ( Y=>nx6210, A=>nx8555);
   i8_r6_lat_q_11_u1 : latchr port map ( QB=>nx8558, D=>nx4356, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(91), A=>nx8558
   );
   i8_r6_lat_q_11_u3 : buf02 port map ( Y=>nx6213, A=>nx8558);
   i7_r17_lat_q_4_u1 : latchr port map ( QB=>nx8561, D=>nx9326, CLK=>nx4270, 
      R=>DecompressedData1(255));
   i7_r17_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(92), A=>nx8561
   );
   i7_r17_lat_q_4_u3 : buf02 port map ( Y=>nx6217, A=>nx8561);
   i8_r6_lat_q_12_u1 : latchr port map ( QB=>nx8564, D=>nx4380, CLK=>nx9362, 
      R=>DecompressedData1(255));
   i8_r6_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(92), A=>nx8564
   );
   i8_r6_lat_q_12_u3 : buf02 port map ( Y=>nx6219, A=>nx8564);
   i7_r16_lat_q_0_u1 : latchr port map ( QB=>nx8567, D=>nx9282, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(96), A=>nx8567
   );
   i7_r16_lat_q_0_u3 : buf02 port map ( Y=>nx6235, A=>nx8567);
   i8_r7_lat_q_0_u1 : latchr port map ( QB=>nx8570, D=>nx4480, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(96), A=>nx8570);
   i8_r7_lat_q_0_u3 : buf02 port map ( Y=>nx6237, A=>nx8570);
   i7_r16_lat_q_1_u1 : latchr port map ( QB=>nx8573, D=>nx9296, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(97), A=>nx8573
   );
   i7_r16_lat_q_1_u3 : buf02 port map ( Y=>nx6240, A=>nx8573);
   i8_r7_lat_q_1_u1 : latchr port map ( QB=>nx8576, D=>nx4504, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(97), A=>nx8576);
   i8_r7_lat_q_1_u3 : buf02 port map ( Y=>nx6243, A=>nx8576);
   i7_r16_lat_q_2_u1 : latchr port map ( QB=>nx8579, D=>nx9306, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(98), A=>nx8579
   );
   i7_r16_lat_q_2_u3 : buf02 port map ( Y=>nx6247, A=>nx8579);
   i8_r7_lat_q_2_u1 : latchr port map ( QB=>nx8582, D=>nx4528, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(98), A=>nx8582);
   i8_r7_lat_q_2_u3 : buf02 port map ( Y=>nx6249, A=>nx8582);
   i7_r16_lat_q_3_u1 : latchr port map ( QB=>nx8585, D=>nx9316, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(99), A=>nx8585
   );
   i7_r16_lat_q_3_u3 : buf02 port map ( Y=>nx6252, A=>nx8585);
   i8_r7_lat_q_3_u1 : latchr port map ( QB=>nx8588, D=>nx4552, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(99), A=>nx8588);
   i8_r7_lat_q_3_u3 : buf02 port map ( Y=>nx6255, A=>nx8588);
   i7_r16_lat_q_4_u1 : latchr port map ( QB=>nx8591, D=>nx9326, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(100), A=>nx8591
   );
   i7_r16_lat_q_4_u3 : buf02 port map ( Y=>nx6259, A=>nx8591);
   i8_r7_lat_q_4_u1 : latchr port map ( QB=>nx8594, D=>nx4576, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(100), A=>nx8594
   );
   i8_r7_lat_q_4_u3 : buf02 port map ( Y=>nx6261, A=>nx8594);
   i7_r16_lat_q_5_u1 : latchr port map ( QB=>nx8597, D=>nx9332, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(101), A=>nx8597
   );
   i7_r16_lat_q_5_u3 : buf02 port map ( Y=>nx6264, A=>nx8597);
   i8_r7_lat_q_5_u1 : latchr port map ( QB=>nx8600, D=>nx4600, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(101), A=>nx8600
   );
   i8_r7_lat_q_5_u3 : buf02 port map ( Y=>nx6267, A=>nx8600);
   i7_r16_lat_q_6_u1 : latchr port map ( QB=>nx8603, D=>nx9336, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(102), A=>nx8603
   );
   i7_r16_lat_q_6_u3 : buf02 port map ( Y=>nx6271, A=>nx8603);
   i8_r7_lat_q_6_u1 : latchr port map ( QB=>nx8606, D=>nx4624, CLK=>nx9364, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(102), A=>nx8606
   );
   i8_r7_lat_q_6_u3 : buf02 port map ( Y=>nx6273, A=>nx8606);
   i7_r16_lat_q_7_u1 : latchr port map ( QB=>nx8609, D=>nx9340, CLK=>nx4454, 
      R=>DecompressedData1(255));
   i7_r16_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(103), A=>nx8609
   );
   i7_r16_lat_q_7_u3 : buf02 port map ( Y=>nx6276, A=>nx8609);
   i8_r7_lat_q_7_u1 : latchr port map ( QB=>nx8612, D=>nx4648, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(103), A=>nx8612
   );
   i8_r7_lat_q_7_u3 : buf02 port map ( Y=>nx6279, A=>nx8612);
   i7_r15_lat_q_0_u1 : latchr port map ( QB=>nx8615, D=>nx9282, CLK=>nx4664, 
      R=>DecompressedData1(255));
   i7_r15_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(104), A=>nx8615
   );
   i7_r15_lat_q_0_u3 : buf02 port map ( Y=>nx6283, A=>nx8615);
   i8_r7_lat_q_8_u1 : latchr port map ( QB=>nx8618, D=>nx4678, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(104), A=>nx8618
   );
   i8_r7_lat_q_8_u3 : buf02 port map ( Y=>nx6285, A=>nx8618);
   i7_r15_lat_q_1_u1 : latchr port map ( QB=>nx8621, D=>nx9296, CLK=>nx4664, 
      R=>DecompressedData1(255));
   i7_r15_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(105), A=>nx8621
   );
   i7_r15_lat_q_1_u3 : buf02 port map ( Y=>nx6288, A=>nx8621);
   i8_r7_lat_q_9_u1 : latchr port map ( QB=>nx8624, D=>nx4702, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(105), A=>nx8624
   );
   i8_r7_lat_q_9_u3 : buf02 port map ( Y=>nx6291, A=>nx8624);
   i7_r15_lat_q_2_u1 : latchr port map ( QB=>nx8627, D=>nx9306, CLK=>nx4664, 
      R=>DecompressedData1(255));
   i7_r15_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(106), A=>nx8627
   );
   i7_r15_lat_q_2_u3 : buf02 port map ( Y=>nx6295, A=>nx8627);
   i8_r7_lat_q_10_u1 : latchr port map ( QB=>nx8630, D=>nx4726, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(106), A=>nx8630
   );
   i8_r7_lat_q_10_u3 : buf02 port map ( Y=>nx6297, A=>nx8630);
   i7_r15_lat_q_3_u1 : latchr port map ( QB=>nx8633, D=>nx9316, CLK=>nx4664, 
      R=>DecompressedData1(255));
   i7_r15_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(107), A=>nx8633
   );
   i7_r15_lat_q_3_u3 : buf02 port map ( Y=>nx6300, A=>nx8633);
   i8_r7_lat_q_11_u1 : latchr port map ( QB=>nx8636, D=>nx4750, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(107), A=>nx8636
   );
   i8_r7_lat_q_11_u3 : buf02 port map ( Y=>nx6303, A=>nx8636);
   i7_r15_lat_q_4_u1 : latchr port map ( QB=>nx8639, D=>nx9326, CLK=>nx4664, 
      R=>DecompressedData1(255));
   i7_r15_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(108), A=>nx8639
   );
   i7_r15_lat_q_4_u3 : buf02 port map ( Y=>nx6307, A=>nx8639);
   i8_r7_lat_q_12_u1 : latchr port map ( QB=>nx8642, D=>nx4774, CLK=>nx9366, 
      R=>DecompressedData1(255));
   i8_r7_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(108), A=>nx8642
   );
   i8_r7_lat_q_12_u3 : buf02 port map ( Y=>nx6309, A=>nx8642);
   i7_r14_lat_q_0_u1 : latchr port map ( QB=>nx8645, D=>nx9284, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(112), A=>nx8645
   );
   i7_r14_lat_q_0_u3 : buf02 port map ( Y=>nx6325, A=>nx8645);
   i8_r8_lat_q_0_u1 : latchr port map ( QB=>nx8648, D=>nx4864, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(112), A=>nx8648
   );
   i8_r8_lat_q_0_u3 : buf02 port map ( Y=>nx6327, A=>nx8648);
   i7_r14_lat_q_1_u1 : latchr port map ( QB=>nx8651, D=>nx9298, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(113), A=>nx8651
   );
   i7_r14_lat_q_1_u3 : buf02 port map ( Y=>nx6331, A=>nx8651);
   i8_r8_lat_q_1_u1 : latchr port map ( QB=>nx8654, D=>nx4888, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(113), A=>nx8654
   );
   i8_r8_lat_q_1_u3 : buf02 port map ( Y=>nx6333, A=>nx8654);
   i7_r14_lat_q_2_u1 : latchr port map ( QB=>nx8657, D=>nx9308, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(114), A=>nx8657
   );
   i7_r14_lat_q_2_u3 : buf02 port map ( Y=>nx6336, A=>nx8657);
   i8_r8_lat_q_2_u1 : latchr port map ( QB=>nx8660, D=>nx4912, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(114), A=>nx8660
   );
   i8_r8_lat_q_2_u3 : buf02 port map ( Y=>nx6339, A=>nx8660);
   i7_r14_lat_q_3_u1 : latchr port map ( QB=>nx8663, D=>nx9318, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(115), A=>nx8663
   );
   i7_r14_lat_q_3_u3 : buf02 port map ( Y=>nx6343, A=>nx8663);
   i8_r8_lat_q_3_u1 : latchr port map ( QB=>nx8666, D=>nx4936, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(115), A=>nx8666
   );
   i8_r8_lat_q_3_u3 : buf02 port map ( Y=>nx6345, A=>nx8666);
   i7_r14_lat_q_4_u1 : latchr port map ( QB=>nx8669, D=>nx9328, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(116), A=>nx8669
   );
   i7_r14_lat_q_4_u3 : buf02 port map ( Y=>nx6348, A=>nx8669);
   i8_r8_lat_q_4_u1 : latchr port map ( QB=>nx8672, D=>nx4960, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(116), A=>nx8672
   );
   i8_r8_lat_q_4_u3 : buf02 port map ( Y=>nx6350, A=>nx8672);
   i7_r14_lat_q_5_u1 : latchr port map ( QB=>nx8675, D=>nx9334, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(117), A=>nx8675
   );
   i7_r14_lat_q_5_u3 : buf02 port map ( Y=>nx6353, A=>nx8675);
   i8_r8_lat_q_5_u1 : latchr port map ( QB=>nx8678, D=>nx4984, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(117), A=>nx8678
   );
   i8_r8_lat_q_5_u3 : buf02 port map ( Y=>nx6355, A=>nx8678);
   i7_r14_lat_q_6_u1 : latchr port map ( QB=>nx8681, D=>nx9338, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(118), A=>nx8681
   );
   i7_r14_lat_q_6_u3 : buf02 port map ( Y=>nx6358, A=>nx8681);
   i8_r8_lat_q_6_u1 : latchr port map ( QB=>nx8684, D=>nx5008, CLK=>nx9368, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(118), A=>nx8684
   );
   i8_r8_lat_q_6_u3 : buf02 port map ( Y=>nx6360, A=>nx8684);
   i7_r14_lat_q_7_u1 : latchr port map ( QB=>nx8687, D=>nx9342, CLK=>nx4838, 
      R=>DecompressedData1(255));
   i7_r14_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(119), A=>nx8687
   );
   i7_r14_lat_q_7_u3 : buf02 port map ( Y=>nx6363, A=>nx8687);
   i8_r8_lat_q_7_u1 : latchr port map ( QB=>nx8690, D=>nx5032, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(119), A=>nx8690
   );
   i8_r8_lat_q_7_u3 : buf02 port map ( Y=>nx6365, A=>nx8690);
   i7_r13_lat_q_0_u1 : latchr port map ( QB=>nx8693, D=>nx9284, CLK=>nx5048, 
      R=>DecompressedData1(255));
   i7_r13_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(120), A=>nx8693
   );
   i7_r13_lat_q_0_u3 : buf02 port map ( Y=>nx6368, A=>nx8693);
   i8_r8_lat_q_8_u1 : latchr port map ( QB=>nx8696, D=>nx5062, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(120), A=>nx8696
   );
   i8_r8_lat_q_8_u3 : buf02 port map ( Y=>nx6370, A=>nx8696);
   i7_r13_lat_q_1_u1 : latchr port map ( QB=>nx8699, D=>nx9298, CLK=>nx5048, 
      R=>DecompressedData1(255));
   i7_r13_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(121), A=>nx8699
   );
   i7_r13_lat_q_1_u3 : buf02 port map ( Y=>nx6373, A=>nx8699);
   i8_r8_lat_q_9_u1 : latchr port map ( QB=>nx8702, D=>nx5086, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(121), A=>nx8702
   );
   i8_r8_lat_q_9_u3 : buf02 port map ( Y=>nx6375, A=>nx8702);
   i7_r13_lat_q_2_u1 : latchr port map ( QB=>nx8705, D=>nx9308, CLK=>nx5048, 
      R=>DecompressedData1(255));
   i7_r13_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(122), A=>nx8705
   );
   i7_r13_lat_q_2_u3 : buf02 port map ( Y=>nx6379, A=>nx8705);
   i8_r8_lat_q_10_u1 : latchr port map ( QB=>nx8708, D=>nx5110, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(122), A=>nx8708
   );
   i8_r8_lat_q_10_u3 : buf02 port map ( Y=>nx6381, A=>nx8708);
   i7_r13_lat_q_3_u1 : latchr port map ( QB=>nx8711, D=>nx9318, CLK=>nx5048, 
      R=>DecompressedData1(255));
   i7_r13_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(123), A=>nx8711
   );
   i7_r13_lat_q_3_u3 : buf02 port map ( Y=>nx6384, A=>nx8711);
   i8_r8_lat_q_11_u1 : latchr port map ( QB=>nx8714, D=>nx5134, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(123), A=>nx8714
   );
   i8_r8_lat_q_11_u3 : buf02 port map ( Y=>nx6387, A=>nx8714);
   i7_r13_lat_q_4_u1 : latchr port map ( QB=>nx8717, D=>nx9328, CLK=>nx5048, 
      R=>DecompressedData1(255));
   i7_r13_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(124), A=>nx8717
   );
   i7_r13_lat_q_4_u3 : buf02 port map ( Y=>nx6391, A=>nx8717);
   i8_r8_lat_q_12_u1 : latchr port map ( QB=>nx8720, D=>nx5158, CLK=>nx9370, 
      R=>DecompressedData1(255));
   i8_r8_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(124), A=>nx8720
   );
   i8_r8_lat_q_12_u3 : buf02 port map ( Y=>nx6393, A=>nx8720);
   i7_r12_lat_q_0_u1 : latchr port map ( QB=>nx8723, D=>nx9284, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(128), A=>nx8723
   );
   i7_r12_lat_q_0_u3 : buf02 port map ( Y=>nx6409, A=>nx8723);
   i8_r9_lat_q_0_u1 : latchr port map ( QB=>nx8726, D=>nx5262, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(128), A=>nx8726
   );
   i8_r9_lat_q_0_u3 : buf02 port map ( Y=>nx6411, A=>nx8726);
   i7_r12_lat_q_1_u1 : latchr port map ( QB=>nx8729, D=>nx9298, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(129), A=>nx8729
   );
   i7_r12_lat_q_1_u3 : buf02 port map ( Y=>nx6415, A=>nx8729);
   i8_r9_lat_q_1_u1 : latchr port map ( QB=>nx8732, D=>nx5286, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(129), A=>nx8732
   );
   i8_r9_lat_q_1_u3 : buf02 port map ( Y=>nx6417, A=>nx8732);
   i7_r12_lat_q_2_u1 : latchr port map ( QB=>nx8735, D=>nx9308, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(130), A=>nx8735
   );
   i7_r12_lat_q_2_u3 : buf02 port map ( Y=>nx6421, A=>nx8735);
   i8_r9_lat_q_2_u1 : latchr port map ( QB=>nx8738, D=>nx5310, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(130), A=>nx8738
   );
   i8_r9_lat_q_2_u3 : buf02 port map ( Y=>nx6423, A=>nx8738);
   i7_r12_lat_q_3_u1 : latchr port map ( QB=>nx8741, D=>nx9318, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(131), A=>nx8741
   );
   i7_r12_lat_q_3_u3 : buf02 port map ( Y=>nx6426, A=>nx8741);
   i8_r9_lat_q_3_u1 : latchr port map ( QB=>nx8744, D=>nx5334, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(131), A=>nx8744
   );
   i8_r9_lat_q_3_u3 : buf02 port map ( Y=>nx6429, A=>nx8744);
   i7_r12_lat_q_4_u1 : latchr port map ( QB=>nx8747, D=>nx9328, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(132), A=>nx8747
   );
   i7_r12_lat_q_4_u3 : buf02 port map ( Y=>nx6433, A=>nx8747);
   i8_r9_lat_q_4_u1 : latchr port map ( QB=>nx8750, D=>nx5358, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(132), A=>nx8750
   );
   i8_r9_lat_q_4_u3 : buf02 port map ( Y=>nx6435, A=>nx8750);
   i7_r12_lat_q_5_u1 : latchr port map ( QB=>nx8753, D=>nx9334, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(133), A=>nx8753
   );
   i7_r12_lat_q_5_u3 : buf02 port map ( Y=>nx6438, A=>nx8753);
   i8_r9_lat_q_5_u1 : latchr port map ( QB=>nx8756, D=>nx5382, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(133), A=>nx8756
   );
   i8_r9_lat_q_5_u3 : buf02 port map ( Y=>nx6441, A=>nx8756);
   i7_r12_lat_q_6_u1 : latchr port map ( QB=>nx8759, D=>nx9338, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(134), A=>nx8759
   );
   i7_r12_lat_q_6_u3 : buf02 port map ( Y=>nx6445, A=>nx8759);
   i8_r9_lat_q_6_u1 : latchr port map ( QB=>nx8762, D=>nx5406, CLK=>nx9372, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(134), A=>nx8762
   );
   i8_r9_lat_q_6_u3 : buf02 port map ( Y=>nx6447, A=>nx8762);
   i7_r12_lat_q_7_u1 : latchr port map ( QB=>nx8765, D=>nx9342, CLK=>nx5228, 
      R=>DecompressedData1(255));
   i7_r12_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(135), A=>nx8765
   );
   i7_r12_lat_q_7_u3 : buf02 port map ( Y=>nx6450, A=>nx8765);
   i8_r9_lat_q_7_u1 : latchr port map ( QB=>nx8768, D=>nx5430, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(135), A=>nx8768
   );
   i8_r9_lat_q_7_u3 : buf02 port map ( Y=>nx6453, A=>nx8768);
   i7_r11_lat_q_0_u1 : latchr port map ( QB=>nx8771, D=>nx9284, CLK=>nx5446, 
      R=>DecompressedData1(255));
   i7_r11_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(136), A=>nx8771
   );
   i7_r11_lat_q_0_u3 : buf02 port map ( Y=>nx6457, A=>nx8771);
   i8_r9_lat_q_8_u1 : latchr port map ( QB=>nx8774, D=>nx5460, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(136), A=>nx8774
   );
   i8_r9_lat_q_8_u3 : buf02 port map ( Y=>nx6459, A=>nx8774);
   i7_r11_lat_q_1_u1 : latchr port map ( QB=>nx8777, D=>nx9298, CLK=>nx5446, 
      R=>DecompressedData1(255));
   i7_r11_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(137), A=>nx8777
   );
   i7_r11_lat_q_1_u3 : buf02 port map ( Y=>nx6462, A=>nx8777);
   i8_r9_lat_q_9_u1 : latchr port map ( QB=>nx8780, D=>nx5484, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(137), A=>nx8780
   );
   i8_r9_lat_q_9_u3 : buf02 port map ( Y=>nx6465, A=>nx8780);
   i7_r11_lat_q_2_u1 : latchr port map ( QB=>nx8783, D=>nx9308, CLK=>nx5446, 
      R=>DecompressedData1(255));
   i7_r11_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(138), A=>nx8783
   );
   i7_r11_lat_q_2_u3 : buf02 port map ( Y=>nx6469, A=>nx8783);
   i8_r9_lat_q_10_u1 : latchr port map ( QB=>nx8786, D=>nx5508, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(138), A=>nx8786
   );
   i8_r9_lat_q_10_u3 : buf02 port map ( Y=>nx6471, A=>nx8786);
   i7_r11_lat_q_3_u1 : latchr port map ( QB=>nx8789, D=>nx9318, CLK=>nx5446, 
      R=>DecompressedData1(255));
   i7_r11_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(139), A=>nx8789
   );
   i7_r11_lat_q_3_u3 : buf02 port map ( Y=>nx6474, A=>nx8789);
   i8_r9_lat_q_11_u1 : latchr port map ( QB=>nx8792, D=>nx5532, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(139), A=>nx8792
   );
   i8_r9_lat_q_11_u3 : buf02 port map ( Y=>nx6477, A=>nx8792);
   i7_r11_lat_q_4_u1 : latchr port map ( QB=>nx8795, D=>nx9328, CLK=>nx5446, 
      R=>DecompressedData1(255));
   i7_r11_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(140), A=>nx8795
   );
   i7_r11_lat_q_4_u3 : buf02 port map ( Y=>nx6481, A=>nx8795);
   i8_r9_lat_q_12_u1 : latchr port map ( QB=>nx8798, D=>nx5556, CLK=>nx9374, 
      R=>DecompressedData1(255));
   i8_r9_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(140), A=>nx8798
   );
   i8_r9_lat_q_12_u3 : buf02 port map ( Y=>nx6483, A=>nx8798);
   i7_r10_lat_q_0_u1 : latchr port map ( QB=>nx8801, D=>nx9284, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(144), A=>nx8801
   );
   i7_r10_lat_q_0_u3 : buf02 port map ( Y=>nx6499, A=>nx8801);
   i8_r10_lat_q_0_u1 : latchr port map ( QB=>nx8804, D=>nx5646, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(144), A=>nx8804
   );
   i8_r10_lat_q_0_u3 : buf02 port map ( Y=>nx6501, A=>nx8804);
   i7_r10_lat_q_1_u1 : latchr port map ( QB=>nx8807, D=>nx9298, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(145), A=>nx8807
   );
   i7_r10_lat_q_1_u3 : buf02 port map ( Y=>nx6505, A=>nx8807);
   i8_r10_lat_q_1_u1 : latchr port map ( QB=>nx8810, D=>nx5670, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(145), A=>nx8810
   );
   i8_r10_lat_q_1_u3 : buf02 port map ( Y=>nx6507, A=>nx8810);
   i7_r10_lat_q_2_u1 : latchr port map ( QB=>nx8813, D=>nx9308, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(146), A=>nx8813
   );
   i7_r10_lat_q_2_u3 : buf02 port map ( Y=>nx6510, A=>nx8813);
   i8_r10_lat_q_2_u1 : latchr port map ( QB=>nx8816, D=>nx5694, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(146), A=>nx8816
   );
   i8_r10_lat_q_2_u3 : buf02 port map ( Y=>nx6513, A=>nx8816);
   i7_r10_lat_q_3_u1 : latchr port map ( QB=>nx8819, D=>nx9318, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(147), A=>nx8819
   );
   i7_r10_lat_q_3_u3 : buf02 port map ( Y=>nx6517, A=>nx8819);
   i8_r10_lat_q_3_u1 : latchr port map ( QB=>nx8822, D=>nx5718, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(147), A=>nx8822
   );
   i8_r10_lat_q_3_u3 : buf02 port map ( Y=>nx6519, A=>nx8822);
   i7_r10_lat_q_4_u1 : latchr port map ( QB=>nx8825, D=>nx9328, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(148), A=>nx8825
   );
   i7_r10_lat_q_4_u3 : buf02 port map ( Y=>nx6522, A=>nx8825);
   i8_r10_lat_q_4_u1 : latchr port map ( QB=>nx8828, D=>nx5742, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(148), A=>nx8828
   );
   i8_r10_lat_q_4_u3 : buf02 port map ( Y=>nx6525, A=>nx8828);
   i7_r10_lat_q_5_u1 : latchr port map ( QB=>nx8831, D=>nx9334, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(149), A=>nx8831
   );
   i7_r10_lat_q_5_u3 : buf02 port map ( Y=>nx6529, A=>nx8831);
   i8_r10_lat_q_5_u1 : latchr port map ( QB=>nx8834, D=>nx5766, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(149), A=>nx8834
   );
   i8_r10_lat_q_5_u3 : buf02 port map ( Y=>nx6531, A=>nx8834);
   i7_r10_lat_q_6_u1 : latchr port map ( QB=>nx8837, D=>nx9338, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(150), A=>nx8837
   );
   i7_r10_lat_q_6_u3 : buf02 port map ( Y=>nx6534, A=>nx8837);
   i8_r10_lat_q_6_u1 : latchr port map ( QB=>nx8840, D=>nx5790, CLK=>nx9376, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(150), A=>nx8840
   );
   i8_r10_lat_q_6_u3 : buf02 port map ( Y=>nx6537, A=>nx8840);
   i7_r10_lat_q_7_u1 : latchr port map ( QB=>nx8843, D=>nx9342, CLK=>nx5620, 
      R=>DecompressedData1(255));
   i7_r10_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(151), A=>nx8843
   );
   i7_r10_lat_q_7_u3 : buf02 port map ( Y=>nx6541, A=>nx8843);
   i8_r10_lat_q_7_u1 : latchr port map ( QB=>nx8846, D=>nx5814, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(151), A=>nx8846
   );
   i8_r10_lat_q_7_u3 : buf02 port map ( Y=>nx6543, A=>nx8846);
   i7_r9_lat_q_0_u1 : latchr port map ( QB=>nx8849, D=>nx9284, CLK=>nx5830, 
      R=>DecompressedData1(255));
   i7_r9_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(152), A=>nx8849
   );
   i7_r9_lat_q_0_u3 : buf02 port map ( Y=>nx6546, A=>nx8849);
   i8_r10_lat_q_8_u1 : latchr port map ( QB=>nx8852, D=>nx5844, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(152), A=>nx8852
   );
   i8_r10_lat_q_8_u3 : buf02 port map ( Y=>nx6549, A=>nx8852);
   i7_r9_lat_q_1_u1 : latchr port map ( QB=>nx8855, D=>nx9298, CLK=>nx5830, 
      R=>DecompressedData1(255));
   i7_r9_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(153), A=>nx8855
   );
   i7_r9_lat_q_1_u3 : buf02 port map ( Y=>nx6553, A=>nx8855);
   i8_r10_lat_q_9_u1 : latchr port map ( QB=>nx8858, D=>nx5868, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(153), A=>nx8858
   );
   i8_r10_lat_q_9_u3 : buf02 port map ( Y=>nx6555, A=>nx8858);
   i7_r9_lat_q_2_u1 : latchr port map ( QB=>nx8861, D=>nx9308, CLK=>nx5830, 
      R=>DecompressedData1(255));
   i7_r9_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(154), A=>nx8861
   );
   i7_r9_lat_q_2_u3 : buf02 port map ( Y=>nx6558, A=>nx8861);
   i8_r10_lat_q_10_u1 : latchr port map ( QB=>nx8864, D=>nx5892, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(154), A=>
      nx8864);
   i8_r10_lat_q_10_u3 : buf02 port map ( Y=>nx6561, A=>nx8864);
   i7_r9_lat_q_3_u1 : latchr port map ( QB=>nx8867, D=>nx9318, CLK=>nx5830, 
      R=>DecompressedData1(255));
   i7_r9_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(155), A=>nx8867
   );
   i7_r9_lat_q_3_u3 : buf02 port map ( Y=>nx6565, A=>nx8867);
   i8_r10_lat_q_11_u1 : latchr port map ( QB=>nx8870, D=>nx5916, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(155), A=>
      nx8870);
   i8_r10_lat_q_11_u3 : buf02 port map ( Y=>nx6567, A=>nx8870);
   i7_r9_lat_q_4_u1 : latchr port map ( QB=>nx8873, D=>nx9328, CLK=>nx5830, 
      R=>DecompressedData1(255));
   i7_r9_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(156), A=>nx8873
   );
   i7_r9_lat_q_4_u3 : buf02 port map ( Y=>nx6570, A=>nx8873);
   i8_r10_lat_q_12_u1 : latchr port map ( QB=>nx8876, D=>nx5940, CLK=>nx9378, 
      R=>DecompressedData1(255));
   i8_r10_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(156), A=>
      nx8876);
   i8_r10_lat_q_12_u3 : buf02 port map ( Y=>nx6573, A=>nx8876);
   i7_r8_lat_q_0_u1 : latchr port map ( QB=>nx8879, D=>nx9284, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(160), A=>nx8879
   );
   i7_r8_lat_q_0_u3 : buf02 port map ( Y=>nx6589, A=>nx8879);
   i8_r11_lat_q_0_u1 : latchr port map ( QB=>nx8882, D=>nx6036, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(160), A=>nx8882
   );
   i8_r11_lat_q_0_u3 : buf02 port map ( Y=>nx6591, A=>nx8882);
   i7_r8_lat_q_1_u1 : latchr port map ( QB=>nx8885, D=>nx9298, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(161), A=>nx8885
   );
   i7_r8_lat_q_1_u3 : buf02 port map ( Y=>nx6594, A=>nx8885);
   i8_r11_lat_q_1_u1 : latchr port map ( QB=>nx8888, D=>nx6060, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(161), A=>nx8888
   );
   i8_r11_lat_q_1_u3 : buf02 port map ( Y=>nx6597, A=>nx8888);
   i7_r8_lat_q_2_u1 : latchr port map ( QB=>nx8891, D=>nx9308, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(162), A=>nx8891
   );
   i7_r8_lat_q_2_u3 : buf02 port map ( Y=>nx6601, A=>nx8891);
   i8_r11_lat_q_2_u1 : latchr port map ( QB=>nx8894, D=>nx6084, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(162), A=>nx8894
   );
   i8_r11_lat_q_2_u3 : buf02 port map ( Y=>nx6603, A=>nx8894);
   i7_r8_lat_q_3_u1 : latchr port map ( QB=>nx8897, D=>nx9318, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(163), A=>nx8897
   );
   i7_r8_lat_q_3_u3 : buf02 port map ( Y=>nx6607, A=>nx8897);
   i8_r11_lat_q_3_u1 : latchr port map ( QB=>nx8900, D=>nx6108, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(163), A=>nx8900
   );
   i8_r11_lat_q_3_u3 : buf02 port map ( Y=>nx6609, A=>nx8900);
   i7_r8_lat_q_4_u1 : latchr port map ( QB=>nx8903, D=>nx9328, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(164), A=>nx8903
   );
   i7_r8_lat_q_4_u3 : buf02 port map ( Y=>nx6612, A=>nx8903);
   i8_r11_lat_q_4_u1 : latchr port map ( QB=>nx8906, D=>nx6132, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(164), A=>nx8906
   );
   i8_r11_lat_q_4_u3 : buf02 port map ( Y=>nx6615, A=>nx8906);
   i7_r8_lat_q_5_u1 : latchr port map ( QB=>nx8909, D=>nx9334, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(165), A=>nx8909
   );
   i7_r8_lat_q_5_u3 : buf02 port map ( Y=>nx6619, A=>nx8909);
   i8_r11_lat_q_5_u1 : latchr port map ( QB=>nx8912, D=>nx6156, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(165), A=>nx8912
   );
   i8_r11_lat_q_5_u3 : buf02 port map ( Y=>nx6621, A=>nx8912);
   i7_r8_lat_q_6_u1 : latchr port map ( QB=>nx8915, D=>nx9338, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(166), A=>nx8915
   );
   i7_r8_lat_q_6_u3 : buf02 port map ( Y=>nx6624, A=>nx8915);
   i8_r11_lat_q_6_u1 : latchr port map ( QB=>nx8918, D=>nx6180, CLK=>nx9380, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(166), A=>nx8918
   );
   i8_r11_lat_q_6_u3 : buf02 port map ( Y=>nx6627, A=>nx8918);
   i7_r8_lat_q_7_u1 : latchr port map ( QB=>nx8921, D=>nx9342, CLK=>nx6010, 
      R=>DecompressedData1(255));
   i7_r8_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(167), A=>nx8921
   );
   i7_r8_lat_q_7_u3 : buf02 port map ( Y=>nx6631, A=>nx8921);
   i8_r11_lat_q_7_u1 : latchr port map ( QB=>nx8924, D=>nx6204, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(167), A=>nx8924
   );
   i8_r11_lat_q_7_u3 : buf02 port map ( Y=>nx6633, A=>nx8924);
   i7_r7_lat_q_0_u1 : latchr port map ( QB=>nx8927, D=>nx9286, CLK=>nx6220, 
      R=>DecompressedData1(255));
   i7_r7_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(168), A=>nx8927
   );
   i7_r7_lat_q_0_u3 : buf02 port map ( Y=>nx6636, A=>nx8927);
   i8_r11_lat_q_8_u1 : latchr port map ( QB=>nx8930, D=>nx6234, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(168), A=>nx8930
   );
   i8_r11_lat_q_8_u3 : buf02 port map ( Y=>nx6639, A=>nx8930);
   i7_r7_lat_q_1_u1 : latchr port map ( QB=>nx8933, D=>nx9300, CLK=>nx6220, 
      R=>DecompressedData1(255));
   i7_r7_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(169), A=>nx8933
   );
   i7_r7_lat_q_1_u3 : buf02 port map ( Y=>nx6643, A=>nx8933);
   i8_r11_lat_q_9_u1 : latchr port map ( QB=>nx8936, D=>nx6258, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(169), A=>nx8936
   );
   i8_r11_lat_q_9_u3 : buf02 port map ( Y=>nx6645, A=>nx8936);
   i7_r7_lat_q_2_u1 : latchr port map ( QB=>nx8939, D=>nx9310, CLK=>nx6220, 
      R=>DecompressedData1(255));
   i7_r7_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(170), A=>nx8939
   );
   i7_r7_lat_q_2_u3 : buf02 port map ( Y=>nx6648, A=>nx8939);
   i8_r11_lat_q_10_u1 : latchr port map ( QB=>nx8942, D=>nx6282, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(170), A=>
      nx8942);
   i8_r11_lat_q_10_u3 : buf02 port map ( Y=>nx6651, A=>nx8942);
   i7_r7_lat_q_3_u1 : latchr port map ( QB=>nx8945, D=>nx9320, CLK=>nx6220, 
      R=>DecompressedData1(255));
   i7_r7_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(171), A=>nx8945
   );
   i7_r7_lat_q_3_u3 : buf02 port map ( Y=>nx6655, A=>nx8945);
   i8_r11_lat_q_11_u1 : latchr port map ( QB=>nx8948, D=>nx6306, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(171), A=>
      nx8948);
   i8_r11_lat_q_11_u3 : buf02 port map ( Y=>nx6657, A=>nx8948);
   i7_r7_lat_q_4_u1 : latchr port map ( QB=>nx8951, D=>nx9330, CLK=>nx6220, 
      R=>DecompressedData1(255));
   i7_r7_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(172), A=>nx8951
   );
   i7_r7_lat_q_4_u3 : buf02 port map ( Y=>nx6660, A=>nx8951);
   i8_r11_lat_q_12_u1 : latchr port map ( QB=>nx8954, D=>nx6330, CLK=>nx9382, 
      R=>DecompressedData1(255));
   i8_r11_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(172), A=>
      nx8954);
   i8_r11_lat_q_12_u3 : buf02 port map ( Y=>nx6663, A=>nx8954);
   i7_r6_lat_q_0_u1 : latchr port map ( QB=>nx8957, D=>nx9286, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(176), A=>nx8957
   );
   i7_r6_lat_q_0_u3 : buf02 port map ( Y=>nx6679, A=>nx8957);
   i8_r12_lat_q_0_u1 : latchr port map ( QB=>nx8960, D=>nx6420, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(176), A=>nx8960
   );
   i8_r12_lat_q_0_u3 : buf02 port map ( Y=>nx6681, A=>nx8960);
   i7_r6_lat_q_1_u1 : latchr port map ( QB=>nx8963, D=>nx9300, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(177), A=>nx8963
   );
   i7_r6_lat_q_1_u3 : buf02 port map ( Y=>nx6684, A=>nx8963);
   i8_r12_lat_q_1_u1 : latchr port map ( QB=>nx8966, D=>nx6444, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(177), A=>nx8966
   );
   i8_r12_lat_q_1_u3 : buf02 port map ( Y=>nx6687, A=>nx8966);
   i7_r6_lat_q_2_u1 : latchr port map ( QB=>nx8969, D=>nx9310, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(178), A=>nx8969
   );
   i7_r6_lat_q_2_u3 : buf02 port map ( Y=>nx6691, A=>nx8969);
   i8_r12_lat_q_2_u1 : latchr port map ( QB=>nx8972, D=>nx6468, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(178), A=>nx8972
   );
   i8_r12_lat_q_2_u3 : buf02 port map ( Y=>nx6693, A=>nx8972);
   i7_r6_lat_q_3_u1 : latchr port map ( QB=>nx8975, D=>nx9320, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(179), A=>nx8975
   );
   i7_r6_lat_q_3_u3 : buf02 port map ( Y=>nx6696, A=>nx8975);
   i8_r12_lat_q_3_u1 : latchr port map ( QB=>nx8978, D=>nx6492, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(179), A=>nx8978
   );
   i8_r12_lat_q_3_u3 : buf02 port map ( Y=>nx6699, A=>nx8978);
   i7_r6_lat_q_4_u1 : latchr port map ( QB=>nx8981, D=>nx9330, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(180), A=>nx8981
   );
   i7_r6_lat_q_4_u3 : buf02 port map ( Y=>nx6703, A=>nx8981);
   i8_r12_lat_q_4_u1 : latchr port map ( QB=>nx8984, D=>nx6516, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(180), A=>nx8984
   );
   i8_r12_lat_q_4_u3 : buf02 port map ( Y=>nx6705, A=>nx8984);
   i7_r6_lat_q_5_u1 : latchr port map ( QB=>nx8987, D=>nx9334, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(181), A=>nx8987
   );
   i7_r6_lat_q_5_u3 : buf02 port map ( Y=>nx6708, A=>nx8987);
   i8_r12_lat_q_5_u1 : latchr port map ( QB=>nx8990, D=>nx6540, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(181), A=>nx8990
   );
   i8_r12_lat_q_5_u3 : buf02 port map ( Y=>nx6711, A=>nx8990);
   i7_r6_lat_q_6_u1 : latchr port map ( QB=>nx8993, D=>nx9338, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(182), A=>nx8993
   );
   i7_r6_lat_q_6_u3 : buf02 port map ( Y=>nx6715, A=>nx8993);
   i8_r12_lat_q_6_u1 : latchr port map ( QB=>nx8996, D=>nx6564, CLK=>nx9384, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(182), A=>nx8996
   );
   i8_r12_lat_q_6_u3 : buf02 port map ( Y=>nx6717, A=>nx8996);
   i7_r6_lat_q_7_u1 : latchr port map ( QB=>nx8999, D=>nx9342, CLK=>nx6394, 
      R=>DecompressedData1(255));
   i7_r6_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(183), A=>nx8999
   );
   i7_r6_lat_q_7_u3 : buf02 port map ( Y=>nx6720, A=>nx8999);
   i8_r12_lat_q_7_u1 : latchr port map ( QB=>nx9002, D=>nx6588, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(183), A=>nx9002
   );
   i8_r12_lat_q_7_u3 : buf02 port map ( Y=>nx6723, A=>nx9002);
   i7_r5_lat_q_0_u1 : latchr port map ( QB=>nx9005, D=>nx9286, CLK=>nx6604, 
      R=>DecompressedData1(255));
   i7_r5_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(184), A=>nx9005
   );
   i7_r5_lat_q_0_u3 : buf02 port map ( Y=>nx6727, A=>nx9005);
   i8_r12_lat_q_8_u1 : latchr port map ( QB=>nx9008, D=>nx6618, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(184), A=>nx9008
   );
   i8_r12_lat_q_8_u3 : buf02 port map ( Y=>nx6729, A=>nx9008);
   i7_r5_lat_q_1_u1 : latchr port map ( QB=>nx9011, D=>nx9300, CLK=>nx6604, 
      R=>DecompressedData1(255));
   i7_r5_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(185), A=>nx9011
   );
   i7_r5_lat_q_1_u3 : buf02 port map ( Y=>nx6732, A=>nx9011);
   i8_r12_lat_q_9_u1 : latchr port map ( QB=>nx9014, D=>nx6642, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(185), A=>nx9014
   );
   i8_r12_lat_q_9_u3 : buf02 port map ( Y=>nx6734, A=>nx9014);
   i7_r5_lat_q_2_u1 : latchr port map ( QB=>nx9017, D=>nx9310, CLK=>nx6604, 
      R=>DecompressedData1(255));
   i7_r5_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(186), A=>nx9017
   );
   i7_r5_lat_q_2_u3 : buf02 port map ( Y=>nx6737, A=>nx9017);
   i8_r12_lat_q_10_u1 : latchr port map ( QB=>nx9020, D=>nx6666, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(186), A=>
      nx9020);
   i8_r12_lat_q_10_u3 : buf02 port map ( Y=>nx6739, A=>nx9020);
   i7_r5_lat_q_3_u1 : latchr port map ( QB=>nx9023, D=>nx9320, CLK=>nx6604, 
      R=>DecompressedData1(255));
   i7_r5_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(187), A=>nx9023
   );
   i7_r5_lat_q_3_u3 : buf02 port map ( Y=>nx6742, A=>nx9023);
   i8_r12_lat_q_11_u1 : latchr port map ( QB=>nx9026, D=>nx6690, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(187), A=>
      nx9026);
   i8_r12_lat_q_11_u3 : buf02 port map ( Y=>nx6744, A=>nx9026);
   i7_r5_lat_q_4_u1 : latchr port map ( QB=>nx9029, D=>nx9330, CLK=>nx6604, 
      R=>DecompressedData1(255));
   i7_r5_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(188), A=>nx9029
   );
   i7_r5_lat_q_4_u3 : buf02 port map ( Y=>nx6747, A=>nx9029);
   i8_r12_lat_q_12_u1 : latchr port map ( QB=>nx9032, D=>nx6714, CLK=>nx9386, 
      R=>DecompressedData1(255));
   i8_r12_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(188), A=>
      nx9032);
   i8_r12_lat_q_12_u3 : buf02 port map ( Y=>nx6749, A=>nx9032);
   i7_r4_lat_q_0_u1 : latchr port map ( QB=>nx9035, D=>nx9286, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(192), A=>nx9035
   );
   i7_r4_lat_q_0_u3 : buf02 port map ( Y=>nx6764, A=>nx9035);
   i8_r13_lat_q_0_u1 : latchr port map ( QB=>nx9038, D=>nx6812, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(192), A=>nx9038
   );
   i8_r13_lat_q_0_u3 : buf02 port map ( Y=>nx6766, A=>nx9038);
   i7_r4_lat_q_1_u1 : latchr port map ( QB=>nx9041, D=>nx9300, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(193), A=>nx9041
   );
   i7_r4_lat_q_1_u3 : buf02 port map ( Y=>nx6769, A=>nx9041);
   i8_r13_lat_q_1_u1 : latchr port map ( QB=>nx9044, D=>nx6836, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(193), A=>nx9044
   );
   i8_r13_lat_q_1_u3 : buf02 port map ( Y=>nx6771, A=>nx9044);
   i7_r4_lat_q_2_u1 : latchr port map ( QB=>nx9047, D=>nx9310, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(194), A=>nx9047
   );
   i7_r4_lat_q_2_u3 : buf02 port map ( Y=>nx6775, A=>nx9047);
   i8_r13_lat_q_2_u1 : latchr port map ( QB=>nx9050, D=>nx6860, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(194), A=>nx9050
   );
   i8_r13_lat_q_2_u3 : buf02 port map ( Y=>nx6777, A=>nx9050);
   i7_r4_lat_q_3_u1 : latchr port map ( QB=>nx9053, D=>nx9320, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(195), A=>nx9053
   );
   i7_r4_lat_q_3_u3 : buf02 port map ( Y=>nx6781, A=>nx9053);
   i8_r13_lat_q_3_u1 : latchr port map ( QB=>nx9056, D=>nx6884, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(195), A=>nx9056
   );
   i8_r13_lat_q_3_u3 : buf02 port map ( Y=>nx6783, A=>nx9056);
   i7_r4_lat_q_4_u1 : latchr port map ( QB=>nx9059, D=>nx9330, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(196), A=>nx9059
   );
   i7_r4_lat_q_4_u3 : buf02 port map ( Y=>nx6787, A=>nx9059);
   i8_r13_lat_q_4_u1 : latchr port map ( QB=>nx9062, D=>nx6908, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(196), A=>nx9062
   );
   i8_r13_lat_q_4_u3 : buf02 port map ( Y=>nx6789, A=>nx9062);
   i7_r4_lat_q_5_u1 : latchr port map ( QB=>nx9065, D=>nx9334, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(197), A=>nx9065
   );
   i7_r4_lat_q_5_u3 : buf02 port map ( Y=>nx6792, A=>nx9065);
   i8_r13_lat_q_5_u1 : latchr port map ( QB=>nx9068, D=>nx6932, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(197), A=>nx9068
   );
   i8_r13_lat_q_5_u3 : buf02 port map ( Y=>nx6794, A=>nx9068);
   i7_r4_lat_q_6_u1 : latchr port map ( QB=>nx9071, D=>nx9338, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(198), A=>nx9071
   );
   i7_r4_lat_q_6_u3 : buf02 port map ( Y=>nx6797, A=>nx9071);
   i8_r13_lat_q_6_u1 : latchr port map ( QB=>nx9074, D=>nx6956, CLK=>nx9388, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(198), A=>nx9074
   );
   i8_r13_lat_q_6_u3 : buf02 port map ( Y=>nx6799, A=>nx9074);
   i7_r4_lat_q_7_u1 : latchr port map ( QB=>nx9077, D=>nx9342, CLK=>nx6786, 
      R=>DecompressedData1(255));
   i7_r4_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(199), A=>nx9077
   );
   i7_r4_lat_q_7_u3 : buf02 port map ( Y=>nx6803, A=>nx9077);
   i8_r13_lat_q_7_u1 : latchr port map ( QB=>nx9080, D=>nx6980, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(199), A=>nx9080
   );
   i8_r13_lat_q_7_u3 : buf02 port map ( Y=>nx6805, A=>nx9080);
   i7_r3_lat_q_0_u1 : latchr port map ( QB=>nx9083, D=>nx9286, CLK=>nx6996, 
      R=>DecompressedData1(255));
   i7_r3_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(200), A=>nx9083
   );
   i7_r3_lat_q_0_u3 : buf02 port map ( Y=>nx6809, A=>nx9083);
   i8_r13_lat_q_8_u1 : latchr port map ( QB=>nx9086, D=>nx7010, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(200), A=>nx9086
   );
   i8_r13_lat_q_8_u3 : buf02 port map ( Y=>nx6811, A=>nx9086);
   i7_r3_lat_q_1_u1 : latchr port map ( QB=>nx9089, D=>nx9300, CLK=>nx6996, 
      R=>DecompressedData1(255));
   i7_r3_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(201), A=>nx9089
   );
   i7_r3_lat_q_1_u3 : buf02 port map ( Y=>nx6815, A=>nx9089);
   i8_r13_lat_q_9_u1 : latchr port map ( QB=>nx9092, D=>nx7034, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(201), A=>nx9092
   );
   i8_r13_lat_q_9_u3 : buf02 port map ( Y=>nx6817, A=>nx9092);
   i7_r3_lat_q_2_u1 : latchr port map ( QB=>nx9095, D=>nx9310, CLK=>nx6996, 
      R=>DecompressedData1(255));
   i7_r3_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(202), A=>nx9095
   );
   i7_r3_lat_q_2_u3 : buf02 port map ( Y=>nx6821, A=>nx9095);
   i8_r13_lat_q_10_u1 : latchr port map ( QB=>nx9098, D=>nx7058, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(202), A=>
      nx9098);
   i8_r13_lat_q_10_u3 : buf02 port map ( Y=>nx6823, A=>nx9098);
   i7_r3_lat_q_3_u1 : latchr port map ( QB=>nx9101, D=>nx9320, CLK=>nx6996, 
      R=>DecompressedData1(255));
   i7_r3_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(203), A=>nx9101
   );
   i7_r3_lat_q_3_u3 : buf02 port map ( Y=>nx6826, A=>nx9101);
   i8_r13_lat_q_11_u1 : latchr port map ( QB=>nx9104, D=>nx7082, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(203), A=>
      nx9104);
   i8_r13_lat_q_11_u3 : buf02 port map ( Y=>nx6828, A=>nx9104);
   i7_r3_lat_q_4_u1 : latchr port map ( QB=>nx9107, D=>nx9330, CLK=>nx6996, 
      R=>DecompressedData1(255));
   i7_r3_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(204), A=>nx9107
   );
   i7_r3_lat_q_4_u3 : buf02 port map ( Y=>nx6831, A=>nx9107);
   i8_r13_lat_q_12_u1 : latchr port map ( QB=>nx9110, D=>nx7106, CLK=>nx9390, 
      R=>DecompressedData1(255));
   i8_r13_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(204), A=>
      nx9110);
   i8_r13_lat_q_12_u3 : buf02 port map ( Y=>nx6833, A=>nx9110);
   i7_r2_lat_q_0_u1 : latchr port map ( QB=>nx9113, D=>nx9286, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(208), A=>nx9113
   );
   i7_r2_lat_q_0_u3 : buf02 port map ( Y=>nx6849, A=>nx9113);
   i8_r14_lat_q_0_u1 : latchr port map ( QB=>nx9116, D=>nx7196, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(208), A=>nx9116
   );
   i8_r14_lat_q_0_u3 : buf02 port map ( Y=>nx6851, A=>nx9116);
   i7_r2_lat_q_1_u1 : latchr port map ( QB=>nx9119, D=>nx9300, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(209), A=>nx9119
   );
   i7_r2_lat_q_1_u3 : buf02 port map ( Y=>nx6854, A=>nx9119);
   i8_r14_lat_q_1_u1 : latchr port map ( QB=>nx9122, D=>nx7220, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(209), A=>nx9122
   );
   i8_r14_lat_q_1_u3 : buf02 port map ( Y=>nx6857, A=>nx9122);
   i7_r2_lat_q_2_u1 : latchr port map ( QB=>nx9125, D=>nx9310, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(210), A=>nx9125
   );
   i7_r2_lat_q_2_u3 : buf02 port map ( Y=>nx6861, A=>nx9125);
   i8_r14_lat_q_2_u1 : latchr port map ( QB=>nx9128, D=>nx7244, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(210), A=>nx9128
   );
   i8_r14_lat_q_2_u3 : buf02 port map ( Y=>nx6863, A=>nx9128);
   i7_r2_lat_q_3_u1 : latchr port map ( QB=>nx9131, D=>nx9320, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(211), A=>nx9131
   );
   i7_r2_lat_q_3_u3 : buf02 port map ( Y=>nx6866, A=>nx9131);
   i8_r14_lat_q_3_u1 : latchr port map ( QB=>nx9134, D=>nx7268, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(211), A=>nx9134
   );
   i8_r14_lat_q_3_u3 : buf02 port map ( Y=>nx6869, A=>nx9134);
   i7_r2_lat_q_4_u1 : latchr port map ( QB=>nx9137, D=>nx9330, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(212), A=>nx9137
   );
   i7_r2_lat_q_4_u3 : buf02 port map ( Y=>nx6873, A=>nx9137);
   i8_r14_lat_q_4_u1 : latchr port map ( QB=>nx9140, D=>nx7292, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(212), A=>nx9140
   );
   i8_r14_lat_q_4_u3 : buf02 port map ( Y=>nx6875, A=>nx9140);
   i7_r2_lat_q_5_u1 : latchr port map ( QB=>nx9143, D=>nx9334, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData1(213), A=>nx9143
   );
   i7_r2_lat_q_5_u3 : buf02 port map ( Y=>nx6878, A=>nx9143);
   i8_r14_lat_q_5_u1 : latchr port map ( QB=>nx9146, D=>nx7316, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(213), A=>nx9146
   );
   i8_r14_lat_q_5_u3 : buf02 port map ( Y=>nx6881, A=>nx9146);
   i7_r2_lat_q_6_u1 : latchr port map ( QB=>nx9149, D=>nx9338, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData1(214), A=>nx9149
   );
   i7_r2_lat_q_6_u3 : buf02 port map ( Y=>nx6885, A=>nx9149);
   i8_r14_lat_q_6_u1 : latchr port map ( QB=>nx9152, D=>nx7340, CLK=>nx9392, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(214), A=>nx9152
   );
   i8_r14_lat_q_6_u3 : buf02 port map ( Y=>nx6887, A=>nx9152);
   i7_r2_lat_q_7_u1 : latchr port map ( QB=>nx9155, D=>nx9342, CLK=>nx7170, 
      R=>DecompressedData1(255));
   i7_r2_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData1(215), A=>nx9155
   );
   i7_r2_lat_q_7_u3 : buf02 port map ( Y=>nx6890, A=>nx9155);
   i8_r14_lat_q_7_u1 : latchr port map ( QB=>nx9158, D=>nx7364, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(215), A=>nx9158
   );
   i8_r14_lat_q_7_u3 : buf02 port map ( Y=>nx6893, A=>nx9158);
   i7_r1_lat_q_0_u1 : latchr port map ( QB=>nx9161, D=>nx9286, CLK=>nx7380, 
      R=>DecompressedData1(255));
   i7_r1_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData1(216), A=>nx9161
   );
   i7_r1_lat_q_0_u3 : buf02 port map ( Y=>nx6897, A=>nx9161);
   i8_r14_lat_q_8_u1 : latchr port map ( QB=>nx9164, D=>nx7394, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(216), A=>nx9164
   );
   i8_r14_lat_q_8_u3 : buf02 port map ( Y=>nx6899, A=>nx9164);
   i7_r1_lat_q_1_u1 : latchr port map ( QB=>nx9167, D=>nx9300, CLK=>nx7380, 
      R=>DecompressedData1(255));
   i7_r1_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData1(217), A=>nx9167
   );
   i7_r1_lat_q_1_u3 : buf02 port map ( Y=>nx6902, A=>nx9167);
   i8_r14_lat_q_9_u1 : latchr port map ( QB=>nx9170, D=>nx7418, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(217), A=>nx9170
   );
   i8_r14_lat_q_9_u3 : buf02 port map ( Y=>nx6905, A=>nx9170);
   i7_r1_lat_q_2_u1 : latchr port map ( QB=>nx9173, D=>nx9310, CLK=>nx7380, 
      R=>DecompressedData1(255));
   i7_r1_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData1(218), A=>nx9173
   );
   i7_r1_lat_q_2_u3 : buf02 port map ( Y=>nx6909, A=>nx9173);
   i8_r14_lat_q_10_u1 : latchr port map ( QB=>nx9176, D=>nx7442, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(218), A=>
      nx9176);
   i8_r14_lat_q_10_u3 : buf02 port map ( Y=>nx6911, A=>nx9176);
   i7_r1_lat_q_3_u1 : latchr port map ( QB=>nx9179, D=>nx9320, CLK=>nx7380, 
      R=>DecompressedData1(255));
   i7_r1_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData1(219), A=>nx9179
   );
   i7_r1_lat_q_3_u3 : buf02 port map ( Y=>nx6914, A=>nx9179);
   i8_r14_lat_q_11_u1 : latchr port map ( QB=>nx9182, D=>nx7466, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(219), A=>
      nx9182);
   i8_r14_lat_q_11_u3 : buf02 port map ( Y=>nx6917, A=>nx9182);
   i7_r1_lat_q_4_u1 : latchr port map ( QB=>nx9185, D=>nx9330, CLK=>nx7380, 
      R=>DecompressedData1(255));
   i7_r1_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData1(220), A=>nx9185
   );
   i7_r1_lat_q_4_u3 : buf02 port map ( Y=>nx6921, A=>nx9185);
   i8_r14_lat_q_12_u1 : latchr port map ( QB=>nx9188, D=>nx7490, CLK=>nx9394, 
      R=>DecompressedData1(255));
   i8_r14_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(220), A=>
      nx9188);
   i8_r14_lat_q_12_u3 : buf02 port map ( Y=>nx6923, A=>nx9188);
   i8_r15_lat_q_0_u1 : latchr port map ( QB=>nx9191, D=>nx1192, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(224), A=>nx9191
   );
   i8_r15_lat_q_0_u3 : buf02 port map ( Y=>nx6939, A=>nx9191);
   i8_r15_lat_q_1_u1 : latchr port map ( QB=>nx9194, D=>nx1206, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(225), A=>nx9194
   );
   i8_r15_lat_q_1_u3 : buf02 port map ( Y=>nx6943, A=>nx9194);
   i8_r15_lat_q_2_u1 : latchr port map ( QB=>nx9197, D=>nx1220, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(226), A=>nx9197
   );
   i8_r15_lat_q_2_u3 : buf02 port map ( Y=>nx6946, A=>nx9197);
   i8_r15_lat_q_3_u1 : latchr port map ( QB=>nx9200, D=>nx1234, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(227), A=>nx9200
   );
   i8_r15_lat_q_3_u3 : buf02 port map ( Y=>nx6949, A=>nx9200);
   i8_r15_lat_q_4_u1 : latchr port map ( QB=>nx9203, D=>nx1248, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(228), A=>nx9203
   );
   i8_r15_lat_q_4_u3 : buf02 port map ( Y=>nx6953, A=>nx9203);
   i8_r15_lat_q_5_u1 : latchr port map ( QB=>nx9206, D=>nx1262, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(229), A=>nx9206
   );
   i8_r15_lat_q_5_u3 : buf02 port map ( Y=>nx6957, A=>nx9206);
   i8_r15_lat_q_6_u1 : latchr port map ( QB=>nx9209, D=>nx1276, CLK=>nx9274, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(230), A=>nx9209
   );
   i8_r15_lat_q_6_u3 : buf02 port map ( Y=>nx6960, A=>nx9209);
   i8_r15_lat_q_7_u1 : latchr port map ( QB=>nx9212, D=>nx1290, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(231), A=>nx9212
   );
   i8_r15_lat_q_7_u3 : buf02 port map ( Y=>nx6963, A=>nx9212);
   i8_r15_lat_q_8_u1 : latchr port map ( QB=>nx9215, D=>nx1304, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(232), A=>nx9215
   );
   i8_r15_lat_q_8_u3 : buf02 port map ( Y=>nx6967, A=>nx9215);
   i8_r15_lat_q_9_u1 : latchr port map ( QB=>nx9218, D=>nx1318, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(233), A=>nx9218
   );
   i8_r15_lat_q_9_u3 : buf02 port map ( Y=>nx6970, A=>nx9218);
   i8_r15_lat_q_10_u1 : latchr port map ( QB=>nx9221, D=>nx1332, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(234), A=>
      nx9221);
   i8_r15_lat_q_10_u3 : buf02 port map ( Y=>nx6973, A=>nx9221);
   i8_r15_lat_q_11_u1 : latchr port map ( QB=>nx9224, D=>nx1346, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(235), A=>
      nx9224);
   i8_r15_lat_q_11_u3 : buf02 port map ( Y=>nx6977, A=>nx9224);
   i8_r15_lat_q_12_u1 : latchr port map ( QB=>nx9227, D=>nx1360, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(236), A=>
      nx9227);
   i8_r15_lat_q_12_u3 : buf02 port map ( Y=>nx6981, A=>nx9227);
   i8_r15_lat_q_13_u1 : latchr port map ( QB=>nx9230, D=>nx1374, CLK=>nx1186, 
      R=>DecompressedData1(255));
   i8_r15_lat_q_13_u2 : inv01 port map ( Y=>DecompressedData2(239), A=>
      nx9230);
   i8_r15_lat_q_13_u3 : buf02 port map ( Y=>nx6984, A=>nx9230);
   i8_r16_lat_q_0_u1 : latchr port map ( QB=>nx9233, D=>nx1398, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_0_u2 : inv01 port map ( Y=>DecompressedData2(240), A=>nx9233
   );
   i8_r16_lat_q_0_u3 : buf02 port map ( Y=>nx6987, A=>nx9233);
   i8_r16_lat_q_1_u1 : latchr port map ( QB=>nx9236, D=>nx1410, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_1_u2 : inv01 port map ( Y=>DecompressedData2(241), A=>nx9236
   );
   i8_r16_lat_q_1_u3 : buf02 port map ( Y=>nx6991, A=>nx9236);
   i8_r16_lat_q_2_u1 : latchr port map ( QB=>nx9239, D=>nx1422, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_2_u2 : inv01 port map ( Y=>DecompressedData2(242), A=>nx9239
   );
   i8_r16_lat_q_2_u3 : buf02 port map ( Y=>nx6995, A=>nx9239);
   i8_r16_lat_q_3_u1 : latchr port map ( QB=>nx9242, D=>nx1434, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_3_u2 : inv01 port map ( Y=>DecompressedData2(243), A=>nx9242
   );
   i8_r16_lat_q_3_u3 : buf02 port map ( Y=>nx6999, A=>nx9242);
   i8_r16_lat_q_4_u1 : latchr port map ( QB=>nx9245, D=>nx1446, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_4_u2 : inv01 port map ( Y=>DecompressedData2(244), A=>nx9245
   );
   i8_r16_lat_q_4_u3 : buf02 port map ( Y=>nx7002, A=>nx9245);
   i8_r16_lat_q_5_u1 : latchr port map ( QB=>nx9248, D=>nx1458, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_5_u2 : inv01 port map ( Y=>DecompressedData2(245), A=>nx9248
   );
   i8_r16_lat_q_5_u3 : buf02 port map ( Y=>nx7005, A=>nx9248);
   i8_r16_lat_q_6_u1 : latchr port map ( QB=>nx9251, D=>nx1470, CLK=>nx9276, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_6_u2 : inv01 port map ( Y=>DecompressedData2(246), A=>nx9251
   );
   i8_r16_lat_q_6_u3 : buf02 port map ( Y=>nx7009, A=>nx9251);
   i8_r16_lat_q_7_u1 : latchr port map ( QB=>nx9254, D=>nx1482, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_7_u2 : inv01 port map ( Y=>DecompressedData2(247), A=>nx9254
   );
   i8_r16_lat_q_7_u3 : buf02 port map ( Y=>nx7013, A=>nx9254);
   i8_r16_lat_q_8_u1 : latchr port map ( QB=>nx9257, D=>nx1494, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_8_u2 : inv01 port map ( Y=>DecompressedData2(248), A=>nx9257
   );
   i8_r16_lat_q_8_u3 : buf02 port map ( Y=>nx7016, A=>nx9257);
   i8_r16_lat_q_9_u1 : latchr port map ( QB=>nx9260, D=>nx1506, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_9_u2 : inv01 port map ( Y=>DecompressedData2(249), A=>nx9260
   );
   i8_r16_lat_q_9_u3 : buf02 port map ( Y=>nx7019, A=>nx9260);
   i8_r16_lat_q_10_u1 : latchr port map ( QB=>nx9263, D=>nx1518, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_10_u2 : inv01 port map ( Y=>DecompressedData2(250), A=>
      nx9263);
   i8_r16_lat_q_10_u3 : buf02 port map ( Y=>nx7023, A=>nx9263);
   i8_r16_lat_q_11_u1 : latchr port map ( QB=>nx9266, D=>nx1530, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_11_u2 : inv01 port map ( Y=>DecompressedData2(251), A=>
      nx9266);
   i8_r16_lat_q_11_u3 : buf02 port map ( Y=>nx7026, A=>nx9266);
   i8_r16_lat_q_12_u1 : latchr port map ( QB=>nx9269, D=>nx1542, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_12_u2 : inv01 port map ( Y=>DecompressedData2(252), A=>
      nx9269);
   i8_r16_lat_q_12_u3 : buf02 port map ( Y=>nx7029, A=>nx9269);
   i8_r16_lat_q_13_u1 : latchr port map ( QB=>nx9272, D=>nx1554, CLK=>nx1394, 
      R=>DecompressedData1(255));
   i8_r16_lat_q_13_u2 : inv01 port map ( Y=>DecompressedData2(255), A=>
      nx9272);
   i8_r16_lat_q_13_u3 : buf02 port map ( Y=>nx7033, A=>nx9272);
   ix9273 : nand02 port map ( Y=>nx9274, A0=>nx5212, A1=>nx5215);
   ix9275 : nand02 port map ( Y=>nx9276, A0=>nx5266, A1=>nx5259);
   ix9277 : inv01 port map ( Y=>nx9278, A=>nx2086);
   ix9279 : inv02 port map ( Y=>nx9280, A=>nx9278);
   ix9281 : inv02 port map ( Y=>nx9282, A=>nx9278);
   ix9283 : inv02 port map ( Y=>nx9284, A=>nx9278);
   ix9285 : inv02 port map ( Y=>nx9286, A=>nx9278);
   ix9287 : inv02 port map ( Y=>nx9288, A=>nx7539);
   ix9289 : inv02 port map ( Y=>nx9290, A=>nx7539);
   ix9291 : inv01 port map ( Y=>nx9292, A=>nx2134);
   ix9293 : inv02 port map ( Y=>nx9294, A=>nx9292);
   ix9295 : inv02 port map ( Y=>nx9296, A=>nx9292);
   ix9297 : inv02 port map ( Y=>nx9298, A=>nx9292);
   ix9299 : inv02 port map ( Y=>nx9300, A=>nx9292);
   ix9301 : inv01 port map ( Y=>nx9302, A=>nx2160);
   ix9303 : inv02 port map ( Y=>nx9304, A=>nx9302);
   ix9305 : inv02 port map ( Y=>nx9306, A=>nx9302);
   ix9307 : inv02 port map ( Y=>nx9308, A=>nx9302);
   ix9309 : inv02 port map ( Y=>nx9310, A=>nx9302);
   ix9311 : inv01 port map ( Y=>nx9312, A=>nx2186);
   ix9313 : inv02 port map ( Y=>nx9314, A=>nx9312);
   ix9315 : inv02 port map ( Y=>nx9316, A=>nx9312);
   ix9317 : inv02 port map ( Y=>nx9318, A=>nx9312);
   ix9319 : inv02 port map ( Y=>nx9320, A=>nx9312);
   ix9321 : inv01 port map ( Y=>nx9322, A=>nx2212);
   ix9323 : inv02 port map ( Y=>nx9324, A=>nx9322);
   ix9325 : inv02 port map ( Y=>nx9326, A=>nx9322);
   ix9327 : inv02 port map ( Y=>nx9328, A=>nx9322);
   ix9329 : inv02 port map ( Y=>nx9330, A=>nx9322);
   ix9331 : inv02 port map ( Y=>nx9332, A=>nx7551);
   ix9333 : inv02 port map ( Y=>nx9334, A=>nx7551);
   ix9335 : inv02 port map ( Y=>nx9336, A=>nx7557);
   ix9337 : inv02 port map ( Y=>nx9338, A=>nx7557);
   ix9339 : inv02 port map ( Y=>nx9340, A=>nx7563);
   ix9341 : inv02 port map ( Y=>nx9342, A=>nx7563);
   ix9343 : inv02 port map ( Y=>nx9344, A=>nx7577);
   ix9345 : inv02 port map ( Y=>nx9346, A=>nx7577);
   ix9347 : inv02 port map ( Y=>nx9348, A=>nx7589);
   ix9349 : inv02 port map ( Y=>nx9350, A=>nx7589);
   ix9351 : inv02 port map ( Y=>nx9352, A=>nx7601);
   ix9353 : inv02 port map ( Y=>nx9354, A=>nx7601);
   ix9355 : inv02 port map ( Y=>nx9356, A=>nx7613);
   ix9357 : inv02 port map ( Y=>nx9358, A=>nx7613);
   ix9359 : inv02 port map ( Y=>nx9360, A=>nx7625);
   ix9361 : inv02 port map ( Y=>nx9362, A=>nx7625);
   ix9363 : inv02 port map ( Y=>nx9364, A=>nx7645);
   ix9365 : inv02 port map ( Y=>nx9366, A=>nx7645);
   ix9367 : inv02 port map ( Y=>nx9368, A=>nx7657);
   ix9369 : inv02 port map ( Y=>nx9370, A=>nx7657);
   ix9371 : inv02 port map ( Y=>nx9372, A=>nx7669);
   ix9373 : inv02 port map ( Y=>nx9374, A=>nx7669);
   ix9375 : inv02 port map ( Y=>nx9376, A=>nx7681);
   ix9377 : inv02 port map ( Y=>nx9378, A=>nx7681);
   ix9379 : inv02 port map ( Y=>nx9380, A=>nx7693);
   ix9381 : inv02 port map ( Y=>nx9382, A=>nx7693);
   ix9383 : inv02 port map ( Y=>nx9384, A=>nx7705);
   ix9385 : inv02 port map ( Y=>nx9386, A=>nx7705);
   ix9387 : inv02 port map ( Y=>nx9388, A=>nx7717);
   ix9389 : inv02 port map ( Y=>nx9390, A=>nx7717);
   ix9391 : inv02 port map ( Y=>nx9392, A=>nx7729);
   ix9393 : inv02 port map ( Y=>nx9394, A=>nx7729);
   ix9395 : inv02 port map ( Y=>nx9396, A=>nx7401);
   ix9397 : inv02 port map ( Y=>nx9398, A=>nx7889);
   ix9399 : inv02 port map ( Y=>nx9400, A=>nx7889);
   ix9401 : inv02 port map ( Y=>nx9402, A=>nx7889);
   ix9403 : inv02 port map ( Y=>nx9404, A=>nx7889);
   ix9405 : inv02 port map ( Y=>nx9406, A=>nx7889);
   ix9407 : inv02 port map ( Y=>nx9408, A=>nx7889);
end arch ;

